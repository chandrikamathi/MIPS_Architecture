
module instruction_mem ( clk, pc, instruction );
  input [7:0] pc;
  output [15:0] instruction;
  input clk;
  wire   n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n4, n5,
         n6, n8, n10, n11, n12, n13, n14;

  INVX2 U3 ( .A(n20), .Y(instruction[5]) );
  OAI21X1 U18 ( .A(n17), .B(n5), .C(n18), .Y(instruction[9]) );
  NAND2X1 U19 ( .A(n19), .B(n20), .Y(instruction[8]) );
  OAI21X1 U20 ( .A(n12), .B(n21), .C(n22), .Y(instruction[7]) );
  NOR2X1 U21 ( .A(instruction[0]), .B(instruction[4]), .Y(n22) );
  OAI21X1 U22 ( .A(n5), .B(n23), .C(n24), .Y(instruction[6]) );
  NOR2X1 U23 ( .A(instruction[1]), .B(instruction[0]), .Y(n24) );
  NAND2X1 U24 ( .A(n25), .B(n12), .Y(n17) );
  NAND2X1 U25 ( .A(n26), .B(n12), .Y(n23) );
  OAI21X1 U26 ( .A(n10), .B(n12), .C(n21), .Y(instruction[3]) );
  OAI21X1 U27 ( .A(pc[1]), .B(n10), .C(n27), .Y(instruction[15]) );
  AOI21X1 U28 ( .A(pc[0]), .B(n25), .C(n4), .Y(n27) );
  NAND3X1 U29 ( .A(n5), .B(n13), .C(n28), .Y(n18) );
  OAI21X1 U30 ( .A(pc[1]), .B(n29), .C(n10), .Y(n28) );
  NOR2X1 U31 ( .A(n5), .B(n20), .Y(instruction[14]) );
  NAND2X1 U32 ( .A(pc[1]), .B(n25), .Y(n20) );
  NOR2X1 U33 ( .A(n13), .B(n10), .Y(n25) );
  OAI21X1 U34 ( .A(n8), .B(n30), .C(n21), .Y(instruction[12]) );
  NAND2X1 U35 ( .A(n5), .B(n12), .Y(n30) );
  OAI21X1 U36 ( .A(n29), .B(pc[2]), .C(n10), .Y(n31) );
  OAI21X1 U37 ( .A(pc[2]), .B(n6), .C(n32), .Y(instruction[11]) );
  NOR2X1 U38 ( .A(instruction[0]), .B(instruction[13]), .Y(n32) );
  NAND3X1 U39 ( .A(n34), .B(n14), .C(n35), .Y(n33) );
  NOR2X1 U40 ( .A(n29), .B(n13), .Y(n35) );
  NOR2X1 U41 ( .A(n34), .B(n10), .Y(instruction[4]) );
  NAND2X1 U42 ( .A(pc[1]), .B(pc[0]), .Y(n34) );
  OAI21X1 U43 ( .A(n12), .B(n36), .C(n37), .Y(instruction[10]) );
  AOI21X1 U44 ( .A(n38), .B(n11), .C(instruction[0]), .Y(n37) );
  NAND3X1 U45 ( .A(n39), .B(n5), .C(n40), .Y(n19) );
  NOR2X1 U46 ( .A(n29), .B(n14), .Y(n40) );
  NOR2X1 U47 ( .A(pc[2]), .B(pc[1]), .Y(n39) );
  NAND2X1 U48 ( .A(n26), .B(n13), .Y(n21) );
  NOR2X1 U49 ( .A(pc[1]), .B(n5), .Y(n38) );
  NAND2X1 U50 ( .A(n26), .B(n5), .Y(n36) );
  NOR2X1 U51 ( .A(n29), .B(pc[3]), .Y(n26) );
  NAND2X1 U52 ( .A(n41), .B(n42), .Y(n29) );
  NOR2X1 U53 ( .A(pc[7]), .B(pc[6]), .Y(n42) );
  NOR2X1 U54 ( .A(pc[5]), .B(pc[4]), .Y(n41) );
  INVX1 U2 ( .A(1'b1), .Y(instruction[2]) );
  INVX2 U5 ( .A(n19), .Y(instruction[0]) );
  INVX2 U6 ( .A(n18), .Y(n4) );
  INVX2 U7 ( .A(pc[0]), .Y(n5) );
  INVX2 U8 ( .A(instruction[4]), .Y(n6) );
  INVX2 U9 ( .A(n33), .Y(instruction[13]) );
  INVX2 U10 ( .A(n31), .Y(n8) );
  INVX2 U11 ( .A(n17), .Y(instruction[1]) );
  INVX2 U12 ( .A(n26), .Y(n10) );
  INVX2 U13 ( .A(n21), .Y(n11) );
  INVX2 U14 ( .A(pc[1]), .Y(n12) );
  INVX2 U15 ( .A(pc[2]), .Y(n13) );
  INVX2 U16 ( .A(pc[3]), .Y(n14) );
endmodule


module IF_stage_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module IF_stage_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:2] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module IF_stage ( clk, rst, instruction_fetch_en, branch_offset_imm, 
        branch_taken, pc, instruction, baseline_en );
  input [5:0] branch_offset_imm;
  output [7:0] pc;
  output [15:0] instruction;
  input clk, rst, instruction_fetch_en, branch_taken;
  output baseline_en;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22,
         N23, N24, n4, n5, n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, n26,
         n28, n30, n32, n34, n36, n38, n39, n7, n9, n11, n13, n15, n17, n19,
         n21, n40, n41, SYNOPSYS_UNCONNECTED_1;

  DFFPOSX1 baseline_en_reg ( .D(n39), .CLK(clk), .Q(baseline_en) );
  DFFSR pc_reg_0_ ( .D(n38), .CLK(clk), .R(n41), .S(1'b1), .Q(pc[0]) );
  DFFSR pc_reg_7_ ( .D(n36), .CLK(clk), .R(n41), .S(1'b1), .Q(pc[7]) );
  DFFSR pc_reg_1_ ( .D(n34), .CLK(clk), .R(n41), .S(1'b1), .Q(pc[1]) );
  DFFSR pc_reg_2_ ( .D(n32), .CLK(clk), .R(n41), .S(1'b1), .Q(pc[2]) );
  DFFSR pc_reg_3_ ( .D(n30), .CLK(clk), .R(n41), .S(1'b1), .Q(pc[3]) );
  DFFSR pc_reg_4_ ( .D(n28), .CLK(clk), .R(n41), .S(1'b1), .Q(pc[4]) );
  DFFSR pc_reg_5_ ( .D(n26), .CLK(clk), .R(n41), .S(1'b1), .Q(pc[5]) );
  DFFSR pc_reg_6_ ( .D(n24), .CLK(clk), .R(n41), .S(1'b1), .Q(pc[6]) );
  OAI21X1 U3 ( .A(instruction_fetch_en), .B(n40), .C(n4), .Y(n24) );
  AOI22X1 U4 ( .A(N23), .B(n5), .C(N15), .D(n6), .Y(n4) );
  OAI21X1 U7 ( .A(instruction_fetch_en), .B(n21), .C(n8), .Y(n26) );
  AOI22X1 U8 ( .A(N22), .B(n5), .C(N14), .D(n6), .Y(n8) );
  OAI21X1 U10 ( .A(instruction_fetch_en), .B(n19), .C(n10), .Y(n28) );
  AOI22X1 U11 ( .A(N21), .B(n5), .C(N13), .D(n6), .Y(n10) );
  OAI21X1 U13 ( .A(instruction_fetch_en), .B(n17), .C(n12), .Y(n30) );
  AOI22X1 U14 ( .A(N20), .B(n5), .C(N12), .D(n6), .Y(n12) );
  OAI21X1 U16 ( .A(instruction_fetch_en), .B(n15), .C(n14), .Y(n32) );
  AOI22X1 U17 ( .A(N19), .B(n5), .C(N11), .D(n6), .Y(n14) );
  OAI21X1 U19 ( .A(instruction_fetch_en), .B(n13), .C(n16), .Y(n34) );
  AOI22X1 U20 ( .A(N18), .B(n5), .C(N10), .D(n6), .Y(n16) );
  OAI21X1 U22 ( .A(instruction_fetch_en), .B(n11), .C(n18), .Y(n36) );
  AOI22X1 U23 ( .A(N24), .B(n5), .C(N16), .D(n6), .Y(n18) );
  OAI21X1 U25 ( .A(instruction_fetch_en), .B(n9), .C(n20), .Y(n38) );
  AOI22X1 U26 ( .A(N17), .B(n5), .C(N9), .D(n6), .Y(n20) );
  AND2X1 U27 ( .A(branch_taken), .B(instruction_fetch_en), .Y(n6) );
  NOR2X1 U28 ( .A(n7), .B(branch_taken), .Y(n5) );
  OAI21X1 U30 ( .A(rst), .B(n7), .C(n22), .Y(n39) );
  NAND2X1 U31 ( .A(baseline_en), .B(rst), .Y(n22) );
  instruction_mem imem ( .clk(clk), .pc(pc), .instruction({instruction[15:3], 
        SYNOPSYS_UNCONNECTED_1, instruction[1:0]}) );
  IF_stage_DW01_inc_0 add_45 ( .A(pc), .SUM({N24, N23, N22, N21, N20, N19, N18, 
        N17}) );
  IF_stage_DW01_add_0 add_42 ( .A(pc), .B({branch_offset_imm[5], 
        branch_offset_imm[5], branch_offset_imm}), .CI(1'b0), .SUM({N16, N15, 
        N14, N13, N12, N11, N10, N9}), .CO() );
  INVX1 U6 ( .A(1'b1), .Y(instruction[2]) );
  INVX2 U12 ( .A(instruction_fetch_en), .Y(n7) );
  INVX2 U18 ( .A(pc[0]), .Y(n9) );
  INVX2 U21 ( .A(pc[7]), .Y(n11) );
  INVX2 U24 ( .A(pc[1]), .Y(n13) );
  INVX2 U29 ( .A(pc[2]), .Y(n15) );
  INVX2 U32 ( .A(pc[3]), .Y(n17) );
  INVX2 U33 ( .A(pc[4]), .Y(n19) );
  INVX2 U42 ( .A(pc[5]), .Y(n21) );
  INVX2 U43 ( .A(pc[6]), .Y(n40) );
  INVX2 U44 ( .A(rst), .Y(n41) );
endmodule


module ID_stage ( clk, rst, baseline_en, pipeline_reg_out, instruction, 
        branch_offset_imm, branch_taken, reg_read_addr_1, reg_read_addr_2, 
        reg_read_data_1, reg_read_data_2 );
  output [57:0] pipeline_reg_out;
  input [15:0] instruction;
  output [5:0] branch_offset_imm;
  output [2:0] reg_read_addr_1;
  output [2:0] reg_read_addr_2;
  input [15:0] reg_read_data_1;
  input [15:0] reg_read_data_2;
  input clk, rst, baseline_en;
  output branch_taken;
  wire   N148, N149, N150, N151, N152, N169, N170, N171, N172, N173, N174,
         N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185,
         N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196,
         N197, N198, N199, N200, N201, N202, N203, N204, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n173, n174;
  wire   [15:9] instruction_reg;

  DFFSR instruction_reg_reg_15_ ( .D(instruction[15]), .CLK(clk), .R(n174), 
        .S(1'b1), .Q(instruction_reg[15]) );
  DFFSR instruction_reg_reg_14_ ( .D(instruction[14]), .CLK(clk), .R(n174), 
        .S(1'b1), .Q(instruction_reg[14]) );
  DFFSR instruction_reg_reg_13_ ( .D(instruction[13]), .CLK(clk), .R(n174), 
        .S(1'b1), .Q(instruction_reg[13]) );
  DFFSR instruction_reg_reg_12_ ( .D(instruction[12]), .CLK(clk), .R(n174), 
        .S(1'b1), .Q(instruction_reg[12]) );
  DFFSR instruction_reg_reg_11_ ( .D(instruction[11]), .CLK(clk), .R(n174), 
        .S(1'b1), .Q(instruction_reg[11]) );
  DFFSR instruction_reg_reg_10_ ( .D(instruction[10]), .CLK(clk), .R(n174), 
        .S(1'b1), .Q(instruction_reg[10]) );
  DFFSR instruction_reg_reg_9_ ( .D(instruction[9]), .CLK(clk), .R(n174), .S(
        1'b1), .Q(instruction_reg[9]) );
  DFFSR instruction_reg_reg_8_ ( .D(instruction[8]), .CLK(clk), .R(n174), .S(
        1'b1), .Q(reg_read_addr_1[2]) );
  DFFSR instruction_reg_reg_7_ ( .D(instruction[7]), .CLK(clk), .R(n174), .S(
        1'b1), .Q(reg_read_addr_1[1]) );
  DFFSR instruction_reg_reg_6_ ( .D(instruction[6]), .CLK(clk), .R(n174), .S(
        1'b1), .Q(reg_read_addr_1[0]) );
  DFFSR instruction_reg_reg_5_ ( .D(instruction[5]), .CLK(clk), .R(n76), .S(
        1'b1), .Q(branch_offset_imm[5]) );
  DFFSR instruction_reg_reg_4_ ( .D(instruction[4]), .CLK(clk), .R(n75), .S(
        1'b1), .Q(branch_offset_imm[4]) );
  DFFSR instruction_reg_reg_3_ ( .D(instruction[3]), .CLK(clk), .R(n174), .S(
        1'b1), .Q(branch_offset_imm[3]) );
  DFFSR instruction_reg_reg_2_ ( .D(instruction[2]), .CLK(clk), .R(n75), .S(
        1'b1), .Q(branch_offset_imm[2]) );
  DFFSR instruction_reg_reg_1_ ( .D(instruction[1]), .CLK(clk), .R(n75), .S(
        1'b1), .Q(branch_offset_imm[1]) );
  DFFSR instruction_reg_reg_0_ ( .D(instruction[0]), .CLK(clk), .R(n174), .S(
        1'b1), .Q(branch_offset_imm[0]) );
  DFFSR pipeline_reg_out_reg_57_ ( .D(baseline_en), .CLK(clk), .R(n174), .S(
        1'b1), .Q(pipeline_reg_out[57]) );
  DFFSR pipeline_reg_out_reg_56_ ( .D(N204), .CLK(clk), .R(n174), .S(1'b1), 
        .Q(pipeline_reg_out[56]) );
  DFFSR pipeline_reg_out_reg_55_ ( .D(N203), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[55]) );
  DFFSR pipeline_reg_out_reg_54_ ( .D(N202), .CLK(clk), .R(n75), .S(1'b1), .Q(
        pipeline_reg_out[54]) );
  DFFSR pipeline_reg_out_reg_53_ ( .D(N201), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[53]) );
  DFFSR pipeline_reg_out_reg_52_ ( .D(N200), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[52]) );
  DFFSR pipeline_reg_out_reg_51_ ( .D(N199), .CLK(clk), .R(n75), .S(1'b1), .Q(
        pipeline_reg_out[51]) );
  DFFSR pipeline_reg_out_reg_50_ ( .D(N198), .CLK(clk), .R(n174), .S(1'b1), 
        .Q(pipeline_reg_out[50]) );
  DFFSR pipeline_reg_out_reg_49_ ( .D(N197), .CLK(clk), .R(n174), .S(1'b1), 
        .Q(pipeline_reg_out[49]) );
  DFFSR pipeline_reg_out_reg_48_ ( .D(N196), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[48]) );
  DFFSR pipeline_reg_out_reg_47_ ( .D(N195), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[47]) );
  DFFSR pipeline_reg_out_reg_46_ ( .D(N194), .CLK(clk), .R(n75), .S(1'b1), .Q(
        pipeline_reg_out[46]) );
  DFFSR pipeline_reg_out_reg_45_ ( .D(N193), .CLK(clk), .R(n174), .S(1'b1), 
        .Q(pipeline_reg_out[45]) );
  DFFSR pipeline_reg_out_reg_44_ ( .D(N192), .CLK(clk), .R(n75), .S(1'b1), .Q(
        pipeline_reg_out[44]) );
  DFFSR pipeline_reg_out_reg_43_ ( .D(N191), .CLK(clk), .R(n174), .S(1'b1), 
        .Q(pipeline_reg_out[43]) );
  DFFSR pipeline_reg_out_reg_42_ ( .D(N190), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[42]) );
  DFFSR pipeline_reg_out_reg_41_ ( .D(N189), .CLK(clk), .R(n174), .S(1'b1), 
        .Q(pipeline_reg_out[41]) );
  DFFSR pipeline_reg_out_reg_40_ ( .D(N188), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[40]) );
  DFFSR pipeline_reg_out_reg_39_ ( .D(N187), .CLK(clk), .R(n174), .S(1'b1), 
        .Q(pipeline_reg_out[39]) );
  DFFSR pipeline_reg_out_reg_38_ ( .D(N186), .CLK(clk), .R(n75), .S(1'b1), .Q(
        pipeline_reg_out[38]) );
  DFFSR pipeline_reg_out_reg_37_ ( .D(N185), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[37]) );
  DFFSR pipeline_reg_out_reg_36_ ( .D(N184), .CLK(clk), .R(n75), .S(1'b1), .Q(
        pipeline_reg_out[36]) );
  DFFSR pipeline_reg_out_reg_35_ ( .D(N183), .CLK(clk), .R(n75), .S(1'b1), .Q(
        pipeline_reg_out[35]) );
  DFFSR pipeline_reg_out_reg_34_ ( .D(N182), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[34]) );
  DFFSR pipeline_reg_out_reg_33_ ( .D(N181), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[33]) );
  DFFSR pipeline_reg_out_reg_32_ ( .D(N180), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[32]) );
  DFFSR pipeline_reg_out_reg_31_ ( .D(N179), .CLK(clk), .R(n174), .S(1'b1), 
        .Q(pipeline_reg_out[31]) );
  DFFSR pipeline_reg_out_reg_30_ ( .D(N178), .CLK(clk), .R(n75), .S(1'b1), .Q(
        pipeline_reg_out[30]) );
  DFFSR pipeline_reg_out_reg_29_ ( .D(N177), .CLK(clk), .R(n174), .S(1'b1), 
        .Q(pipeline_reg_out[29]) );
  DFFSR pipeline_reg_out_reg_28_ ( .D(N176), .CLK(clk), .R(n75), .S(1'b1), .Q(
        pipeline_reg_out[28]) );
  DFFSR pipeline_reg_out_reg_27_ ( .D(N175), .CLK(clk), .R(n174), .S(1'b1), 
        .Q(pipeline_reg_out[27]) );
  DFFSR pipeline_reg_out_reg_26_ ( .D(N174), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[26]) );
  DFFSR pipeline_reg_out_reg_25_ ( .D(N173), .CLK(clk), .R(n75), .S(1'b1), .Q(
        pipeline_reg_out[25]) );
  DFFSR pipeline_reg_out_reg_24_ ( .D(N172), .CLK(clk), .R(n174), .S(1'b1), 
        .Q(pipeline_reg_out[24]) );
  DFFSR pipeline_reg_out_reg_23_ ( .D(N171), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[23]) );
  DFFSR pipeline_reg_out_reg_22_ ( .D(N170), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[22]) );
  DFFSR pipeline_reg_out_reg_21_ ( .D(N169), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[21]) );
  DFFSR pipeline_reg_out_reg_20_ ( .D(n78), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[20]) );
  DFFSR pipeline_reg_out_reg_19_ ( .D(n79), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[19]) );
  DFFSR pipeline_reg_out_reg_18_ ( .D(n81), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[18]) );
  DFFSR pipeline_reg_out_reg_17_ ( .D(n83), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[17]) );
  DFFSR pipeline_reg_out_reg_16_ ( .D(n85), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[16]) );
  DFFSR pipeline_reg_out_reg_15_ ( .D(n87), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[15]) );
  DFFSR pipeline_reg_out_reg_14_ ( .D(n89), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[14]) );
  DFFSR pipeline_reg_out_reg_13_ ( .D(n91), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[13]) );
  DFFSR pipeline_reg_out_reg_12_ ( .D(n93), .CLK(clk), .R(n76), .S(1'b1), .Q(
        pipeline_reg_out[12]) );
  DFFSR pipeline_reg_out_reg_11_ ( .D(n95), .CLK(clk), .R(n75), .S(1'b1), .Q(
        pipeline_reg_out[11]) );
  DFFSR pipeline_reg_out_reg_10_ ( .D(n97), .CLK(clk), .R(n75), .S(1'b1), .Q(
        pipeline_reg_out[10]) );
  DFFSR pipeline_reg_out_reg_9_ ( .D(n99), .CLK(clk), .R(n75), .S(1'b1), .Q(
        pipeline_reg_out[9]) );
  DFFSR pipeline_reg_out_reg_8_ ( .D(n101), .CLK(clk), .R(n75), .S(1'b1), .Q(
        pipeline_reg_out[8]) );
  DFFSR pipeline_reg_out_reg_7_ ( .D(n103), .CLK(clk), .R(n75), .S(1'b1), .Q(
        pipeline_reg_out[7]) );
  DFFSR pipeline_reg_out_reg_6_ ( .D(n104), .CLK(clk), .R(n75), .S(1'b1), .Q(
        pipeline_reg_out[6]) );
  DFFSR pipeline_reg_out_reg_5_ ( .D(n106), .CLK(clk), .R(n75), .S(1'b1), .Q(
        pipeline_reg_out[5]) );
  DFFSR pipeline_reg_out_reg_4_ ( .D(N152), .CLK(clk), .R(n75), .S(1'b1), .Q(
        pipeline_reg_out[4]) );
  DFFSR pipeline_reg_out_reg_3_ ( .D(N151), .CLK(clk), .R(n75), .S(1'b1), .Q(
        pipeline_reg_out[3]) );
  DFFSR pipeline_reg_out_reg_2_ ( .D(N150), .CLK(clk), .R(n75), .S(1'b1), .Q(
        pipeline_reg_out[2]) );
  DFFSR pipeline_reg_out_reg_1_ ( .D(N149), .CLK(clk), .R(n75), .S(1'b1), .Q(
        pipeline_reg_out[1]) );
  DFFSR pipeline_reg_out_reg_0_ ( .D(N148), .CLK(clk), .R(n75), .S(1'b1), .Q(
        pipeline_reg_out[0]) );
  OR2X2 U77 ( .A(n138), .B(n107), .Y(n172) );
  OAI22X1 U123 ( .A(n110), .B(n118), .C(n120), .D(n115), .Y(reg_read_addr_2[2]) );
  OAI22X1 U124 ( .A(n110), .B(n119), .C(n120), .D(n116), .Y(reg_read_addr_2[1]) );
  OAI22X1 U125 ( .A(n110), .B(n173), .C(n120), .D(n117), .Y(reg_read_addr_2[0]) );
  NOR2X1 U126 ( .A(n121), .B(n122), .Y(branch_taken) );
  NAND3X1 U127 ( .A(n123), .B(n124), .C(n125), .Y(n122) );
  NOR2X1 U128 ( .A(n126), .B(n127), .Y(n125) );
  NAND2X1 U129 ( .A(n105), .B(n86), .Y(n127) );
  NAND3X1 U130 ( .A(n82), .B(n80), .C(n84), .Y(n126) );
  NOR2X1 U131 ( .A(instruction_reg[10]), .B(n128), .Y(n124) );
  NAND2X1 U132 ( .A(n115), .B(n117), .Y(n128) );
  NOR2X1 U133 ( .A(n107), .B(n129), .Y(n123) );
  NAND3X1 U134 ( .A(n130), .B(n131), .C(n132), .Y(n121) );
  NOR2X1 U135 ( .A(n133), .B(n134), .Y(n132) );
  NAND3X1 U136 ( .A(n96), .B(n94), .C(n98), .Y(n134) );
  NAND3X1 U137 ( .A(n90), .B(n88), .C(n92), .Y(n133) );
  NOR2X1 U138 ( .A(reg_read_data_1[1]), .B(n135), .Y(n131) );
  NAND2X1 U139 ( .A(n102), .B(n100), .Y(n135) );
  NOR2X1 U140 ( .A(reg_read_data_1[15]), .B(reg_read_data_1[14]), .Y(n130) );
  AOI21X1 U141 ( .A(n136), .B(n137), .C(n138), .Y(N204) );
  NAND3X1 U142 ( .A(n139), .B(n107), .C(instruction_reg[14]), .Y(n137) );
  AOI21X1 U143 ( .A(n136), .B(n140), .C(n138), .Y(N203) );
  NAND2X1 U144 ( .A(n141), .B(n107), .Y(n140) );
  OAI21X1 U145 ( .A(n114), .B(n113), .C(n129), .Y(n141) );
  AOI21X1 U146 ( .A(n136), .B(n142), .C(n138), .Y(N202) );
  OAI21X1 U147 ( .A(instruction_reg[13]), .B(instruction_reg[14]), .C(n143), 
        .Y(n142) );
  NOR2X1 U148 ( .A(instruction_reg[15]), .B(instruction_reg[12]), .Y(n143) );
  NAND3X1 U149 ( .A(instruction_reg[15]), .B(n111), .C(n112), .Y(n136) );
  AND2X1 U150 ( .A(baseline_en), .B(reg_read_data_1[15]), .Y(N201) );
  AND2X1 U151 ( .A(baseline_en), .B(reg_read_data_1[14]), .Y(N200) );
  NOR2X1 U152 ( .A(n77), .B(n80), .Y(N199) );
  NOR2X1 U153 ( .A(n77), .B(n82), .Y(N198) );
  NOR2X1 U154 ( .A(n77), .B(n84), .Y(N197) );
  NOR2X1 U155 ( .A(n77), .B(n86), .Y(N196) );
  NOR2X1 U156 ( .A(n77), .B(n88), .Y(N195) );
  NOR2X1 U157 ( .A(n77), .B(n90), .Y(N194) );
  NOR2X1 U158 ( .A(n77), .B(n92), .Y(N193) );
  NOR2X1 U159 ( .A(n77), .B(n94), .Y(N192) );
  NOR2X1 U160 ( .A(n77), .B(n96), .Y(N191) );
  NOR2X1 U161 ( .A(n77), .B(n98), .Y(N190) );
  NOR2X1 U162 ( .A(n77), .B(n100), .Y(N189) );
  NOR2X1 U163 ( .A(n77), .B(n102), .Y(N188) );
  AND2X1 U164 ( .A(baseline_en), .B(reg_read_data_1[1]), .Y(N187) );
  NOR2X1 U165 ( .A(n77), .B(n105), .Y(N186) );
  OAI21X1 U166 ( .A(n109), .B(n144), .C(n145), .Y(N185) );
  OAI21X1 U167 ( .A(n109), .B(n146), .C(n145), .Y(N184) );
  OAI21X1 U168 ( .A(n109), .B(n147), .C(n145), .Y(N183) );
  OAI21X1 U169 ( .A(n109), .B(n148), .C(n145), .Y(N182) );
  OAI21X1 U170 ( .A(n109), .B(n149), .C(n145), .Y(N181) );
  OAI21X1 U171 ( .A(n109), .B(n150), .C(n145), .Y(N180) );
  OAI21X1 U172 ( .A(n109), .B(n151), .C(n145), .Y(N179) );
  OAI21X1 U173 ( .A(n109), .B(n152), .C(n145), .Y(N178) );
  OAI21X1 U174 ( .A(n109), .B(n153), .C(n145), .Y(N177) );
  OAI21X1 U175 ( .A(n109), .B(n154), .C(n145), .Y(N176) );
  OAI21X1 U176 ( .A(n109), .B(n155), .C(n145), .Y(N175) );
  NAND2X1 U177 ( .A(n108), .B(branch_offset_imm[5]), .Y(n145) );
  OAI22X1 U178 ( .A(n109), .B(n156), .C(n119), .D(n157), .Y(N174) );
  OAI22X1 U179 ( .A(n109), .B(n158), .C(n173), .D(n157), .Y(N173) );
  OAI21X1 U180 ( .A(n109), .B(n159), .C(n160), .Y(N172) );
  NAND2X1 U181 ( .A(branch_offset_imm[2]), .B(n108), .Y(n160) );
  OAI21X1 U182 ( .A(n109), .B(n161), .C(n162), .Y(N171) );
  NAND2X1 U183 ( .A(branch_offset_imm[1]), .B(n108), .Y(n162) );
  OAI21X1 U184 ( .A(n109), .B(n163), .C(n164), .Y(N170) );
  NAND2X1 U185 ( .A(branch_offset_imm[0]), .B(n108), .Y(n164) );
  NAND2X1 U186 ( .A(n109), .B(baseline_en), .Y(n157) );
  NAND3X1 U187 ( .A(n166), .B(n174), .C(instruction_reg[15]), .Y(n165) );
  OAI21X1 U188 ( .A(instruction_reg[14]), .B(n112), .C(n129), .Y(n166) );
  NAND2X1 U189 ( .A(instruction_reg[14]), .B(n112), .Y(n129) );
  NOR2X1 U190 ( .A(n120), .B(n77), .Y(N169) );
  NAND3X1 U191 ( .A(instruction_reg[15]), .B(instruction_reg[13]), .C(n167), 
        .Y(n120) );
  NOR2X1 U192 ( .A(instruction_reg[14]), .B(n114), .Y(n167) );
  NAND2X1 U193 ( .A(reg_read_data_2[15]), .B(baseline_en), .Y(n144) );
  NAND2X1 U194 ( .A(reg_read_data_2[14]), .B(baseline_en), .Y(n146) );
  NAND2X1 U195 ( .A(reg_read_data_2[13]), .B(baseline_en), .Y(n147) );
  NAND2X1 U196 ( .A(reg_read_data_2[12]), .B(baseline_en), .Y(n148) );
  NAND2X1 U197 ( .A(reg_read_data_2[11]), .B(baseline_en), .Y(n149) );
  NAND2X1 U198 ( .A(reg_read_data_2[10]), .B(baseline_en), .Y(n150) );
  NAND2X1 U199 ( .A(reg_read_data_2[9]), .B(baseline_en), .Y(n151) );
  NAND2X1 U200 ( .A(reg_read_data_2[8]), .B(baseline_en), .Y(n152) );
  NAND2X1 U201 ( .A(reg_read_data_2[7]), .B(baseline_en), .Y(n153) );
  NAND2X1 U202 ( .A(reg_read_data_2[6]), .B(baseline_en), .Y(n154) );
  NAND2X1 U203 ( .A(reg_read_data_2[5]), .B(baseline_en), .Y(n155) );
  NAND2X1 U204 ( .A(reg_read_data_2[4]), .B(baseline_en), .Y(n156) );
  NAND2X1 U205 ( .A(reg_read_data_2[3]), .B(baseline_en), .Y(n158) );
  NAND2X1 U206 ( .A(reg_read_data_2[2]), .B(baseline_en), .Y(n159) );
  NAND2X1 U207 ( .A(reg_read_data_2[1]), .B(baseline_en), .Y(n161) );
  NAND2X1 U208 ( .A(reg_read_data_2[0]), .B(baseline_en), .Y(n163) );
  NOR2X1 U209 ( .A(n138), .B(n168), .Y(N152) );
  OAI21X1 U210 ( .A(n169), .B(n107), .C(n170), .Y(n168) );
  NAND3X1 U211 ( .A(n111), .B(n107), .C(n112), .Y(n170) );
  NAND2X1 U212 ( .A(n113), .B(n114), .Y(n139) );
  AOI21X1 U213 ( .A(instruction_reg[13]), .B(instruction_reg[12]), .C(
        instruction_reg[14]), .Y(n169) );
  NOR2X1 U214 ( .A(n115), .B(n77), .Y(N151) );
  NOR2X1 U215 ( .A(n116), .B(n77), .Y(N150) );
  NOR2X1 U216 ( .A(n117), .B(n77), .Y(N149) );
  NOR2X1 U217 ( .A(n171), .B(n172), .Y(N148) );
  NAND2X1 U218 ( .A(baseline_en), .B(n174), .Y(n138) );
  NAND3X1 U219 ( .A(n114), .B(n111), .C(instruction_reg[13]), .Y(n171) );
  BUFX2 U78 ( .A(n174), .Y(n75) );
  BUFX2 U79 ( .A(n174), .Y(n76) );
  INVX2 U80 ( .A(n165), .Y(n109) );
  INVX2 U81 ( .A(baseline_en), .Y(n77) );
  INVX2 U82 ( .A(n144), .Y(n78) );
  INVX2 U83 ( .A(n146), .Y(n79) );
  INVX2 U84 ( .A(reg_read_data_1[13]), .Y(n80) );
  INVX2 U85 ( .A(n147), .Y(n81) );
  INVX2 U86 ( .A(reg_read_data_1[12]), .Y(n82) );
  INVX2 U87 ( .A(n148), .Y(n83) );
  INVX2 U88 ( .A(reg_read_data_1[11]), .Y(n84) );
  INVX2 U89 ( .A(n149), .Y(n85) );
  INVX2 U90 ( .A(reg_read_data_1[10]), .Y(n86) );
  INVX2 U91 ( .A(n150), .Y(n87) );
  INVX2 U92 ( .A(reg_read_data_1[9]), .Y(n88) );
  INVX2 U93 ( .A(n151), .Y(n89) );
  INVX2 U94 ( .A(reg_read_data_1[8]), .Y(n90) );
  INVX2 U95 ( .A(n152), .Y(n91) );
  INVX2 U96 ( .A(reg_read_data_1[7]), .Y(n92) );
  INVX2 U97 ( .A(n153), .Y(n93) );
  INVX2 U98 ( .A(reg_read_data_1[6]), .Y(n94) );
  INVX2 U99 ( .A(n154), .Y(n95) );
  INVX2 U100 ( .A(reg_read_data_1[5]), .Y(n96) );
  INVX2 U101 ( .A(n155), .Y(n97) );
  INVX2 U102 ( .A(reg_read_data_1[4]), .Y(n98) );
  INVX2 U103 ( .A(n156), .Y(n99) );
  INVX2 U104 ( .A(reg_read_data_1[3]), .Y(n100) );
  INVX2 U105 ( .A(n158), .Y(n101) );
  INVX2 U106 ( .A(reg_read_data_1[2]), .Y(n102) );
  INVX2 U107 ( .A(n159), .Y(n103) );
  INVX2 U108 ( .A(n161), .Y(n104) );
  INVX2 U109 ( .A(reg_read_data_1[0]), .Y(n105) );
  INVX2 U110 ( .A(n163), .Y(n106) );
  INVX2 U111 ( .A(instruction_reg[15]), .Y(n107) );
  INVX2 U112 ( .A(n157), .Y(n108) );
  INVX2 U113 ( .A(n120), .Y(n110) );
  INVX2 U114 ( .A(instruction_reg[14]), .Y(n111) );
  INVX2 U115 ( .A(n139), .Y(n112) );
  INVX2 U116 ( .A(instruction_reg[13]), .Y(n113) );
  INVX2 U117 ( .A(instruction_reg[12]), .Y(n114) );
  INVX2 U118 ( .A(instruction_reg[11]), .Y(n115) );
  INVX2 U119 ( .A(instruction_reg[10]), .Y(n116) );
  INVX2 U120 ( .A(instruction_reg[9]), .Y(n117) );
  INVX2 U121 ( .A(branch_offset_imm[5]), .Y(n118) );
  INVX2 U122 ( .A(branch_offset_imm[4]), .Y(n119) );
  INVX2 U220 ( .A(branch_offset_imm[3]), .Y(n173) );
  INVX2 U221 ( .A(rst), .Y(n174) );
endmodule


module alu_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [15:0] A;
  input [15:0] SH;
  output [15:0] B;
  input DATA_TC, SH_TC;
  wire   ML_int_1__0_, ML_int_2__1_, ML_int_2__0_, ML_int_3__3_, ML_int_3__2_,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120;
  wire   [4:0] SHMAG;

  MUX2X1 M1_3_15 ( .B(n1), .A(n25), .S(n49), .Y(n54) );
  MUX2X1 M1_3_14 ( .B(n4), .A(n28), .S(n49), .Y(n55) );
  MUX2X1 M1_3_13 ( .B(n7), .A(n31), .S(n49), .Y(n56) );
  MUX2X1 M1_3_12 ( .B(n10), .A(n34), .S(n49), .Y(n57) );
  MUX2X1 M1_3_11 ( .B(n13), .A(ML_int_3__3_), .S(n49), .Y(n58) );
  MUX2X1 M1_3_10 ( .B(n16), .A(ML_int_3__2_), .S(n49), .Y(n59) );
  MUX2X1 M1_3_9 ( .B(n19), .A(n44), .S(n49), .Y(n60) );
  MUX2X1 M1_3_8 ( .B(n22), .A(n45), .S(n49), .Y(n61) );
  MUX2X1 M1_2_15 ( .B(n2), .A(n14), .S(n48), .Y(n62) );
  MUX2X1 M1_2_14 ( .B(n5), .A(n17), .S(n48), .Y(n63) );
  MUX2X1 M1_2_13 ( .B(n8), .A(n20), .S(n48), .Y(n64) );
  MUX2X1 M1_2_12 ( .B(n11), .A(n23), .S(n48), .Y(n65) );
  MUX2X1 M1_2_11 ( .B(n14), .A(n26), .S(n48), .Y(n66) );
  MUX2X1 M1_2_10 ( .B(n17), .A(n29), .S(n48), .Y(n67) );
  MUX2X1 M1_2_9 ( .B(n20), .A(n32), .S(n48), .Y(n68) );
  MUX2X1 M1_2_8 ( .B(n23), .A(n35), .S(n48), .Y(n69) );
  MUX2X1 M1_2_7 ( .B(n26), .A(n37), .S(n48), .Y(n70) );
  MUX2X1 M1_2_6 ( .B(n29), .A(n40), .S(n48), .Y(n71) );
  MUX2X1 M1_2_5 ( .B(n32), .A(ML_int_2__1_), .S(n48), .Y(n72) );
  MUX2X1 M1_2_4 ( .B(n35), .A(ML_int_2__0_), .S(n48), .Y(n73) );
  MUX2X1 M1_1_15 ( .B(n3), .A(n9), .S(n47), .Y(n74) );
  MUX2X1 M1_1_14 ( .B(n6), .A(n12), .S(n47), .Y(n75) );
  MUX2X1 M1_1_13 ( .B(n9), .A(n15), .S(n47), .Y(n76) );
  MUX2X1 M1_1_12 ( .B(n12), .A(n18), .S(n47), .Y(n77) );
  MUX2X1 M1_1_11 ( .B(n15), .A(n21), .S(n47), .Y(n78) );
  MUX2X1 M1_1_10 ( .B(n18), .A(n24), .S(n47), .Y(n79) );
  MUX2X1 M1_1_9 ( .B(n21), .A(n27), .S(n47), .Y(n80) );
  MUX2X1 M1_1_8 ( .B(n24), .A(n30), .S(n47), .Y(n81) );
  MUX2X1 M1_1_7 ( .B(n27), .A(n33), .S(n47), .Y(n82) );
  MUX2X1 M1_1_6 ( .B(n30), .A(n36), .S(n47), .Y(n83) );
  MUX2X1 M1_1_5 ( .B(n33), .A(n39), .S(n47), .Y(n84) );
  MUX2X1 M1_1_4 ( .B(n36), .A(n42), .S(n47), .Y(n85) );
  MUX2X1 M1_1_3 ( .B(n39), .A(n43), .S(n47), .Y(n86) );
  MUX2X1 M1_1_2 ( .B(n42), .A(ML_int_1__0_), .S(n47), .Y(n87) );
  MUX2X1 M1_0_15 ( .B(A[15]), .A(A[14]), .S(n46), .Y(n88) );
  MUX2X1 M1_0_14 ( .B(A[14]), .A(A[13]), .S(n46), .Y(n89) );
  MUX2X1 M1_0_13 ( .B(A[13]), .A(A[12]), .S(n46), .Y(n90) );
  MUX2X1 M1_0_12 ( .B(A[12]), .A(A[11]), .S(n46), .Y(n91) );
  MUX2X1 M1_0_11 ( .B(A[11]), .A(A[10]), .S(n46), .Y(n92) );
  MUX2X1 M1_0_10 ( .B(A[10]), .A(A[9]), .S(n46), .Y(n93) );
  MUX2X1 M1_0_9 ( .B(A[9]), .A(A[8]), .S(n46), .Y(n94) );
  MUX2X1 M1_0_8 ( .B(A[8]), .A(A[7]), .S(n46), .Y(n95) );
  MUX2X1 M1_0_7 ( .B(A[7]), .A(A[6]), .S(n46), .Y(n96) );
  MUX2X1 M1_0_6 ( .B(A[6]), .A(A[5]), .S(n46), .Y(n97) );
  MUX2X1 M1_0_5 ( .B(A[5]), .A(A[4]), .S(n46), .Y(n98) );
  MUX2X1 M1_0_4 ( .B(A[4]), .A(A[3]), .S(n46), .Y(n99) );
  MUX2X1 M1_0_3 ( .B(A[3]), .A(A[2]), .S(n46), .Y(n100) );
  MUX2X1 M1_0_2 ( .B(A[2]), .A(A[1]), .S(n46), .Y(n101) );
  MUX2X1 M1_0_1 ( .B(A[1]), .A(A[0]), .S(n46), .Y(n102) );
  INVX2 U3 ( .A(SHMAG[0]), .Y(n46) );
  INVX2 U4 ( .A(SHMAG[1]), .Y(n47) );
  INVX2 U5 ( .A(SHMAG[2]), .Y(n48) );
  INVX2 U6 ( .A(SHMAG[3]), .Y(n49) );
  INVX2 U7 ( .A(n62), .Y(n1) );
  INVX2 U8 ( .A(n74), .Y(n2) );
  INVX2 U9 ( .A(n88), .Y(n3) );
  INVX2 U10 ( .A(n63), .Y(n4) );
  INVX2 U11 ( .A(n75), .Y(n5) );
  INVX2 U12 ( .A(n89), .Y(n6) );
  INVX2 U13 ( .A(n64), .Y(n7) );
  INVX2 U14 ( .A(n76), .Y(n8) );
  INVX2 U15 ( .A(n90), .Y(n9) );
  INVX2 U16 ( .A(n65), .Y(n10) );
  INVX2 U17 ( .A(n77), .Y(n11) );
  INVX2 U18 ( .A(n91), .Y(n12) );
  INVX2 U19 ( .A(n66), .Y(n13) );
  INVX2 U20 ( .A(n78), .Y(n14) );
  INVX2 U21 ( .A(n92), .Y(n15) );
  INVX2 U22 ( .A(n67), .Y(n16) );
  INVX2 U23 ( .A(n79), .Y(n17) );
  INVX2 U24 ( .A(n93), .Y(n18) );
  INVX2 U25 ( .A(n68), .Y(n19) );
  INVX2 U26 ( .A(n80), .Y(n20) );
  INVX2 U27 ( .A(n94), .Y(n21) );
  INVX2 U28 ( .A(n69), .Y(n22) );
  INVX2 U29 ( .A(n81), .Y(n23) );
  INVX2 U30 ( .A(n95), .Y(n24) );
  INVX2 U31 ( .A(n70), .Y(n25) );
  INVX2 U32 ( .A(n82), .Y(n26) );
  INVX2 U33 ( .A(n96), .Y(n27) );
  INVX2 U34 ( .A(n71), .Y(n28) );
  INVX2 U35 ( .A(n83), .Y(n29) );
  INVX2 U36 ( .A(n97), .Y(n30) );
  INVX2 U37 ( .A(n72), .Y(n31) );
  INVX2 U38 ( .A(n84), .Y(n32) );
  INVX2 U39 ( .A(n98), .Y(n33) );
  INVX2 U40 ( .A(n73), .Y(n34) );
  INVX2 U41 ( .A(n85), .Y(n35) );
  INVX2 U42 ( .A(n99), .Y(n36) );
  INVX2 U43 ( .A(n86), .Y(n37) );
  INVX2 U44 ( .A(ML_int_3__3_), .Y(n38) );
  INVX2 U45 ( .A(n100), .Y(n39) );
  INVX2 U46 ( .A(n87), .Y(n40) );
  INVX2 U47 ( .A(ML_int_3__2_), .Y(n41) );
  INVX2 U48 ( .A(n101), .Y(n42) );
  INVX2 U49 ( .A(n102), .Y(n43) );
  INVX2 U50 ( .A(n105), .Y(n44) );
  INVX2 U51 ( .A(n106), .Y(n45) );
  INVX2 U52 ( .A(n114), .Y(n50) );
  INVX2 U53 ( .A(SH[15]), .Y(n51) );
  INVX2 U54 ( .A(SH[12]), .Y(n52) );
  INVX2 U55 ( .A(SH[7]), .Y(n53) );
  NOR2X1 U56 ( .A(n60), .B(n103), .Y(B[9]) );
  NOR2X1 U57 ( .A(n61), .B(n103), .Y(B[8]) );
  NOR2X1 U58 ( .A(n70), .B(n104), .Y(B[7]) );
  NOR2X1 U59 ( .A(n71), .B(n104), .Y(B[6]) );
  NOR2X1 U60 ( .A(n72), .B(n104), .Y(B[5]) );
  NOR2X1 U61 ( .A(n73), .B(n104), .Y(B[4]) );
  NOR2X1 U62 ( .A(n104), .B(n38), .Y(B[3]) );
  NOR2X1 U63 ( .A(n104), .B(n41), .Y(B[2]) );
  NOR2X1 U64 ( .A(n104), .B(n105), .Y(B[1]) );
  NOR2X1 U65 ( .A(n54), .B(n103), .Y(B[15]) );
  NOR2X1 U66 ( .A(n55), .B(n103), .Y(B[14]) );
  NOR2X1 U67 ( .A(n56), .B(n103), .Y(B[13]) );
  NOR2X1 U68 ( .A(n57), .B(n103), .Y(B[12]) );
  NOR2X1 U69 ( .A(n58), .B(n103), .Y(B[11]) );
  NOR2X1 U70 ( .A(n59), .B(n103), .Y(B[10]) );
  NOR2X1 U71 ( .A(n104), .B(n106), .Y(B[0]) );
  OR2X1 U72 ( .A(n103), .B(n49), .Y(n104) );
  AOI21X1 U73 ( .A(n107), .B(SH[3]), .C(n50), .Y(SHMAG[3]) );
  NAND2X1 U74 ( .A(SHMAG[4]), .B(n51), .Y(n103) );
  AOI21X1 U75 ( .A(n107), .B(SH[4]), .C(n50), .Y(SHMAG[4]) );
  NOR2X1 U76 ( .A(n48), .B(n86), .Y(ML_int_3__3_) );
  NOR2X1 U77 ( .A(n48), .B(n87), .Y(ML_int_3__2_) );
  NAND2X1 U78 ( .A(ML_int_2__1_), .B(SHMAG[2]), .Y(n105) );
  NAND2X1 U79 ( .A(ML_int_2__0_), .B(SHMAG[2]), .Y(n106) );
  AOI21X1 U80 ( .A(n107), .B(SH[2]), .C(n50), .Y(SHMAG[2]) );
  NOR2X1 U81 ( .A(n47), .B(n102), .Y(ML_int_2__1_) );
  AND2X1 U82 ( .A(ML_int_1__0_), .B(SHMAG[1]), .Y(ML_int_2__0_) );
  AOI21X1 U83 ( .A(n107), .B(SH[1]), .C(n50), .Y(SHMAG[1]) );
  AND2X1 U84 ( .A(A[0]), .B(SHMAG[0]), .Y(ML_int_1__0_) );
  OAI21X1 U85 ( .A(SH[0]), .B(n50), .C(n107), .Y(SHMAG[0]) );
  OAI21X1 U86 ( .A(n108), .B(n109), .C(SH[15]), .Y(n107) );
  NAND3X1 U87 ( .A(SH[9]), .B(SH[8]), .C(n110), .Y(n109) );
  NOR2X1 U88 ( .A(n53), .B(n111), .Y(n110) );
  NAND2X1 U89 ( .A(SH[6]), .B(SH[5]), .Y(n111) );
  NAND3X1 U90 ( .A(SH[14]), .B(SH[13]), .C(n112), .Y(n108) );
  NOR2X1 U91 ( .A(n52), .B(n113), .Y(n112) );
  NAND2X1 U92 ( .A(SH[11]), .B(SH[10]), .Y(n113) );
  OAI21X1 U93 ( .A(n115), .B(n116), .C(n51), .Y(n114) );
  NAND3X1 U94 ( .A(n117), .B(n52), .C(n118), .Y(n116) );
  NOR2X1 U95 ( .A(SH[11]), .B(SH[10]), .Y(n118) );
  NOR2X1 U96 ( .A(SH[14]), .B(SH[13]), .Y(n117) );
  NAND3X1 U97 ( .A(n119), .B(n53), .C(n120), .Y(n115) );
  NOR2X1 U98 ( .A(SH[6]), .B(SH[5]), .Y(n120) );
  NOR2X1 U99 ( .A(SH[9]), .B(SH[8]), .Y(n119) );
endmodule


module alu_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [15:2] carry;

  FAX1 U2_15 ( .A(A[15]), .B(n2), .C(carry[15]), .YC(), .YS(DIFF[15]) );
  FAX1 U2_14 ( .A(A[14]), .B(n3), .C(carry[14]), .YC(carry[15]), .YS(DIFF[14])
         );
  FAX1 U2_13 ( .A(A[13]), .B(n4), .C(carry[13]), .YC(carry[14]), .YS(DIFF[13])
         );
  FAX1 U2_12 ( .A(A[12]), .B(n5), .C(carry[12]), .YC(carry[13]), .YS(DIFF[12])
         );
  FAX1 U2_11 ( .A(A[11]), .B(n6), .C(carry[11]), .YC(carry[12]), .YS(DIFF[11])
         );
  FAX1 U2_10 ( .A(A[10]), .B(n7), .C(carry[10]), .YC(carry[11]), .YS(DIFF[10])
         );
  FAX1 U2_9 ( .A(A[9]), .B(n8), .C(carry[9]), .YC(carry[10]), .YS(DIFF[9]) );
  FAX1 U2_8 ( .A(A[8]), .B(n9), .C(carry[8]), .YC(carry[9]), .YS(DIFF[8]) );
  FAX1 U2_7 ( .A(A[7]), .B(n10), .C(carry[7]), .YC(carry[8]), .YS(DIFF[7]) );
  FAX1 U2_6 ( .A(A[6]), .B(n11), .C(carry[6]), .YC(carry[7]), .YS(DIFF[6]) );
  FAX1 U2_5 ( .A(A[5]), .B(n12), .C(carry[5]), .YC(carry[6]), .YS(DIFF[5]) );
  FAX1 U2_4 ( .A(A[4]), .B(n13), .C(carry[4]), .YC(carry[5]), .YS(DIFF[4]) );
  FAX1 U2_3 ( .A(A[3]), .B(n14), .C(carry[3]), .YC(carry[4]), .YS(DIFF[3]) );
  FAX1 U2_2 ( .A(A[2]), .B(n15), .C(carry[2]), .YC(carry[3]), .YS(DIFF[2]) );
  FAX1 U2_1 ( .A(A[1]), .B(n16), .C(n1), .YC(carry[2]), .YS(DIFF[1]) );
  OR2X2 U1 ( .A(A[0]), .B(n17), .Y(n1) );
  XNOR2X1 U2 ( .A(n17), .B(A[0]), .Y(DIFF[0]) );
  INVX2 U3 ( .A(B[15]), .Y(n2) );
  INVX2 U4 ( .A(B[14]), .Y(n3) );
  INVX2 U5 ( .A(B[13]), .Y(n4) );
  INVX2 U6 ( .A(B[12]), .Y(n5) );
  INVX2 U7 ( .A(B[11]), .Y(n6) );
  INVX2 U8 ( .A(B[10]), .Y(n7) );
  INVX2 U9 ( .A(B[9]), .Y(n8) );
  INVX2 U10 ( .A(B[8]), .Y(n9) );
  INVX2 U11 ( .A(B[7]), .Y(n10) );
  INVX2 U12 ( .A(B[6]), .Y(n11) );
  INVX2 U13 ( .A(B[5]), .Y(n12) );
  INVX2 U14 ( .A(B[4]), .Y(n13) );
  INVX2 U15 ( .A(B[3]), .Y(n14) );
  INVX2 U16 ( .A(B[2]), .Y(n15) );
  INVX2 U17 ( .A(B[1]), .Y(n16) );
  INVX2 U18 ( .A(B[0]), .Y(n17) );
endmodule


module alu_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [15:2] carry;

  FAX1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .YC(), .YS(SUM[15]) );
  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YC(carry[15]), .YS(
        SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module alu ( a, b, cmd, r );
  input [15:0] a;
  input [15:0] b;
  input [2:0] cmd;
  output [15:0] r;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N113, N114, N115, N116, N117, N118, N119, N120,
         N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131,
         N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142,
         N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153,
         N154, N155, N156, N157, N158, N159, N160, n74, n75, n76, n77, n78,
         n79, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n80, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432;

  NAND3X1 U54 ( .A(n74), .B(n75), .C(n76), .Y(r[9]) );
  AOI21X1 U55 ( .A(N42), .B(n322), .C(n311), .Y(n76) );
  AOI22X1 U56 ( .A(N122), .B(n325), .C(N58), .D(n323), .Y(n77) );
  AOI22X1 U57 ( .A(a[9]), .B(n78), .C(b[9]), .D(n79), .Y(n75) );
  OAI21X1 U58 ( .A(n341), .B(n3), .C(n81), .Y(n79) );
  AOI21X1 U59 ( .A(n326), .B(n341), .C(n321), .Y(n81) );
  OAI21X1 U60 ( .A(b[9]), .B(n82), .C(n83), .Y(n78) );
  AOI22X1 U61 ( .A(N154), .B(n328), .C(N138), .D(n327), .Y(n74) );
  NAND3X1 U62 ( .A(n84), .B(n85), .C(n86), .Y(r[8]) );
  AOI21X1 U63 ( .A(N41), .B(n322), .C(n312), .Y(n86) );
  AOI22X1 U64 ( .A(N121), .B(n325), .C(N57), .D(n323), .Y(n87) );
  AOI22X1 U65 ( .A(a[8]), .B(n88), .C(b[8]), .D(n89), .Y(n85) );
  OAI21X1 U66 ( .A(n3), .B(n342), .C(n90), .Y(n89) );
  AOI21X1 U67 ( .A(n326), .B(n342), .C(n321), .Y(n90) );
  OAI21X1 U68 ( .A(b[8]), .B(n82), .C(n83), .Y(n88) );
  AOI22X1 U69 ( .A(N153), .B(n328), .C(N137), .D(n327), .Y(n84) );
  NAND3X1 U70 ( .A(n91), .B(n92), .C(n93), .Y(r[7]) );
  AOI21X1 U71 ( .A(N40), .B(n322), .C(n313), .Y(n93) );
  AOI22X1 U72 ( .A(N120), .B(n325), .C(N56), .D(n323), .Y(n94) );
  AOI22X1 U73 ( .A(n32), .B(n95), .C(b[7]), .D(n96), .Y(n92) );
  OAI21X1 U74 ( .A(n3), .B(n28), .C(n97), .Y(n96) );
  AOI21X1 U75 ( .A(n326), .B(n28), .C(n321), .Y(n97) );
  OAI21X1 U76 ( .A(b[7]), .B(n82), .C(n83), .Y(n95) );
  AOI22X1 U77 ( .A(N152), .B(n328), .C(N136), .D(n327), .Y(n91) );
  NAND3X1 U78 ( .A(n98), .B(n99), .C(n100), .Y(r[6]) );
  AOI21X1 U79 ( .A(N39), .B(n322), .C(n314), .Y(n100) );
  AOI22X1 U80 ( .A(N119), .B(n325), .C(N55), .D(n323), .Y(n101) );
  AOI22X1 U81 ( .A(n27), .B(n102), .C(b[6]), .D(n103), .Y(n99) );
  OAI21X1 U82 ( .A(n3), .B(n26), .C(n104), .Y(n103) );
  AOI21X1 U83 ( .A(n326), .B(n26), .C(n321), .Y(n104) );
  OAI21X1 U84 ( .A(b[6]), .B(n82), .C(n83), .Y(n102) );
  AOI22X1 U85 ( .A(N151), .B(n328), .C(N135), .D(n327), .Y(n98) );
  NAND3X1 U86 ( .A(n105), .B(n106), .C(n107), .Y(r[5]) );
  AOI21X1 U87 ( .A(N38), .B(n322), .C(n315), .Y(n107) );
  AOI22X1 U88 ( .A(N118), .B(n325), .C(N54), .D(n323), .Y(n108) );
  AOI22X1 U89 ( .A(n25), .B(n109), .C(b[5]), .D(n110), .Y(n106) );
  OAI21X1 U90 ( .A(n3), .B(n24), .C(n111), .Y(n110) );
  AOI21X1 U91 ( .A(n326), .B(n24), .C(n321), .Y(n111) );
  OAI21X1 U92 ( .A(b[5]), .B(n82), .C(n83), .Y(n109) );
  AOI22X1 U93 ( .A(N150), .B(n328), .C(N134), .D(n327), .Y(n105) );
  NAND3X1 U94 ( .A(n112), .B(n113), .C(n114), .Y(r[4]) );
  AOI21X1 U95 ( .A(N37), .B(n322), .C(n316), .Y(n114) );
  AOI22X1 U96 ( .A(N117), .B(n325), .C(N53), .D(n323), .Y(n115) );
  AOI22X1 U97 ( .A(a[4]), .B(n116), .C(n15), .D(n117), .Y(n113) );
  OAI21X1 U98 ( .A(n3), .B(n22), .C(n118), .Y(n117) );
  AOI21X1 U99 ( .A(n326), .B(n22), .C(n321), .Y(n118) );
  OAI21X1 U100 ( .A(n15), .B(n82), .C(n83), .Y(n116) );
  AOI22X1 U101 ( .A(N149), .B(n328), .C(N133), .D(n327), .Y(n112) );
  NAND3X1 U102 ( .A(n119), .B(n120), .C(n121), .Y(r[3]) );
  AOI21X1 U103 ( .A(N36), .B(n322), .C(n317), .Y(n121) );
  AOI22X1 U104 ( .A(N116), .B(n325), .C(N52), .D(n323), .Y(n122) );
  AOI22X1 U105 ( .A(n21), .B(n123), .C(n13), .D(n124), .Y(n120) );
  OAI21X1 U106 ( .A(n3), .B(n20), .C(n125), .Y(n124) );
  AOI21X1 U107 ( .A(n326), .B(n20), .C(n321), .Y(n125) );
  OAI21X1 U108 ( .A(n13), .B(n82), .C(n83), .Y(n123) );
  AOI22X1 U109 ( .A(N148), .B(n328), .C(N132), .D(n327), .Y(n119) );
  NAND3X1 U110 ( .A(n126), .B(n127), .C(n128), .Y(r[2]) );
  AOI21X1 U111 ( .A(N35), .B(n322), .C(n318), .Y(n128) );
  AOI22X1 U112 ( .A(N115), .B(n325), .C(N51), .D(n323), .Y(n129) );
  AOI22X1 U113 ( .A(a[2]), .B(n130), .C(n11), .D(n131), .Y(n127) );
  OAI21X1 U114 ( .A(n3), .B(n18), .C(n132), .Y(n131) );
  AOI21X1 U115 ( .A(n326), .B(n18), .C(n321), .Y(n132) );
  OAI21X1 U116 ( .A(n11), .B(n82), .C(n83), .Y(n130) );
  AOI22X1 U117 ( .A(N147), .B(n328), .C(N131), .D(n327), .Y(n126) );
  NAND3X1 U118 ( .A(n133), .B(n134), .C(n135), .Y(r[1]) );
  AOI21X1 U119 ( .A(N34), .B(n322), .C(n319), .Y(n135) );
  AOI22X1 U120 ( .A(N114), .B(n325), .C(N50), .D(n323), .Y(n136) );
  AOI22X1 U121 ( .A(n17), .B(n137), .C(n9), .D(n138), .Y(n134) );
  OAI21X1 U122 ( .A(n3), .B(n16), .C(n139), .Y(n138) );
  AOI21X1 U123 ( .A(n326), .B(n16), .C(n321), .Y(n139) );
  OAI21X1 U124 ( .A(n9), .B(n82), .C(n83), .Y(n137) );
  AOI22X1 U125 ( .A(N146), .B(n328), .C(N130), .D(n327), .Y(n133) );
  NAND3X1 U126 ( .A(n140), .B(n141), .C(n142), .Y(r[15]) );
  AOI21X1 U127 ( .A(N48), .B(n322), .C(n305), .Y(n142) );
  AOI22X1 U128 ( .A(N128), .B(n325), .C(N64), .D(n323), .Y(n143) );
  AOI22X1 U129 ( .A(n34), .B(n144), .C(b[15]), .D(n145), .Y(n141) );
  OAI21X1 U130 ( .A(n3), .B(n33), .C(n146), .Y(n145) );
  AOI21X1 U131 ( .A(n326), .B(n33), .C(n321), .Y(n146) );
  OAI21X1 U132 ( .A(b[15]), .B(n82), .C(n83), .Y(n144) );
  AOI22X1 U133 ( .A(N160), .B(n328), .C(N144), .D(n327), .Y(n140) );
  NAND3X1 U134 ( .A(n147), .B(n148), .C(n149), .Y(r[14]) );
  AOI21X1 U135 ( .A(N47), .B(n322), .C(n306), .Y(n149) );
  AOI22X1 U136 ( .A(N127), .B(n325), .C(N63), .D(n323), .Y(n150) );
  AOI22X1 U137 ( .A(a[14]), .B(n151), .C(b[14]), .D(n152), .Y(n148) );
  OAI21X1 U138 ( .A(n3), .B(n293), .C(n153), .Y(n152) );
  AOI21X1 U139 ( .A(n326), .B(n293), .C(n321), .Y(n153) );
  OAI21X1 U140 ( .A(b[14]), .B(n82), .C(n83), .Y(n151) );
  AOI22X1 U141 ( .A(N159), .B(n328), .C(N143), .D(n327), .Y(n147) );
  NAND3X1 U142 ( .A(n154), .B(n155), .C(n156), .Y(r[13]) );
  AOI21X1 U143 ( .A(N46), .B(n322), .C(n307), .Y(n156) );
  AOI22X1 U144 ( .A(N126), .B(n325), .C(N62), .D(n323), .Y(n157) );
  AOI22X1 U145 ( .A(a[13]), .B(n158), .C(b[13]), .D(n159), .Y(n155) );
  OAI21X1 U146 ( .A(n3), .B(n336), .C(n160), .Y(n159) );
  AOI21X1 U147 ( .A(n326), .B(n336), .C(n321), .Y(n160) );
  OAI21X1 U148 ( .A(b[13]), .B(n82), .C(n83), .Y(n158) );
  AOI22X1 U149 ( .A(N158), .B(n328), .C(N142), .D(n327), .Y(n154) );
  NAND3X1 U150 ( .A(n161), .B(n162), .C(n163), .Y(r[12]) );
  AOI21X1 U151 ( .A(N45), .B(n322), .C(n308), .Y(n163) );
  AOI22X1 U152 ( .A(N125), .B(n325), .C(N61), .D(n323), .Y(n164) );
  AOI22X1 U153 ( .A(a[12]), .B(n165), .C(b[12]), .D(n166), .Y(n162) );
  OAI21X1 U154 ( .A(n3), .B(n289), .C(n167), .Y(n166) );
  AOI21X1 U155 ( .A(n326), .B(n289), .C(n321), .Y(n167) );
  OAI21X1 U156 ( .A(b[12]), .B(n82), .C(n83), .Y(n165) );
  AOI22X1 U157 ( .A(N157), .B(n328), .C(N141), .D(n327), .Y(n161) );
  NAND3X1 U158 ( .A(n168), .B(n169), .C(n170), .Y(r[11]) );
  AOI21X1 U159 ( .A(N44), .B(n322), .C(n309), .Y(n170) );
  AOI22X1 U160 ( .A(N124), .B(n325), .C(N60), .D(n323), .Y(n171) );
  AOI22X1 U161 ( .A(a[11]), .B(n172), .C(b[11]), .D(n173), .Y(n169) );
  OAI21X1 U162 ( .A(n3), .B(n339), .C(n174), .Y(n173) );
  AOI21X1 U163 ( .A(n326), .B(n339), .C(n321), .Y(n174) );
  OAI21X1 U164 ( .A(b[11]), .B(n82), .C(n83), .Y(n172) );
  AOI22X1 U165 ( .A(N156), .B(n328), .C(N140), .D(n327), .Y(n168) );
  NAND3X1 U166 ( .A(n175), .B(n176), .C(n177), .Y(r[10]) );
  AOI21X1 U167 ( .A(N43), .B(n322), .C(n310), .Y(n177) );
  AOI22X1 U168 ( .A(N123), .B(n325), .C(N59), .D(n323), .Y(n178) );
  AOI22X1 U169 ( .A(a[10]), .B(n179), .C(b[10]), .D(n180), .Y(n176) );
  OAI21X1 U170 ( .A(n3), .B(n287), .C(n181), .Y(n180) );
  AOI21X1 U171 ( .A(n326), .B(n287), .C(n321), .Y(n181) );
  OAI21X1 U172 ( .A(b[10]), .B(n82), .C(n83), .Y(n179) );
  AOI22X1 U173 ( .A(N155), .B(n328), .C(N139), .D(n327), .Y(n175) );
  NAND3X1 U174 ( .A(n182), .B(n183), .C(n184), .Y(r[0]) );
  AOI21X1 U175 ( .A(N33), .B(n322), .C(n320), .Y(n184) );
  AOI22X1 U176 ( .A(N113), .B(n325), .C(N49), .D(n323), .Y(n185) );
  NAND3X1 U177 ( .A(n329), .B(n324), .C(cmd[0]), .Y(n186) );
  NAND3X1 U178 ( .A(cmd[2]), .B(n329), .C(cmd[0]), .Y(n187) );
  NAND3X1 U179 ( .A(n329), .B(n324), .C(n330), .Y(n188) );
  AOI22X1 U180 ( .A(a[0]), .B(n189), .C(n7), .D(n190), .Y(n183) );
  OAI21X1 U181 ( .A(n3), .B(n344), .C(n191), .Y(n190) );
  AOI21X1 U182 ( .A(n326), .B(n344), .C(n321), .Y(n191) );
  OAI21X1 U184 ( .A(n7), .B(n82), .C(n83), .Y(n189) );
  NAND3X1 U185 ( .A(cmd[0]), .B(n324), .C(cmd[1]), .Y(n83) );
  NAND3X1 U186 ( .A(n330), .B(n329), .C(cmd[2]), .Y(n82) );
  AOI22X1 U187 ( .A(N145), .B(n328), .C(N129), .D(n327), .Y(n182) );
  NAND3X1 U188 ( .A(cmd[2]), .B(n330), .C(cmd[1]), .Y(n192) );
  NAND3X1 U189 ( .A(cmd[0]), .B(cmd[2]), .C(cmd[1]), .Y(n193) );
  alu_DW01_ash_0 sll_36 ( .A({n34, a[14:8], n32, a[6], n25, n23, n21, n19, n17, 
        a[0]}), .DATA_TC(1'b0), .SH({b[15:5], n15, n13, n11, n9, n7}), .SH_TC(
        1'b0), .B({N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, 
        N118, N117, N116, N115, N114, N113}) );
  alu_DW01_sub_0 sub_28 ( .A({n34, a[14:8], n32, n27, a[5], n23, a[3], n19, 
        n17, a[0]}), .B({b[15:5], n15, n13, n11, n9, n7}), .CI(1'b0), .DIFF({
        N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, 
        N50, N49}), .CO() );
  alu_DW01_add_0 add_26 ( .A({a[15:8], n32, n27, a[5], n23, a[3], n19, n17, 
        a[0]}), .B({b[15:5], n15, n13, n11, n9, n7}), .CI(1'b0), .SUM({N48, 
        N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, 
        N33}), .CO() );
  OR2X2 U2 ( .A(n6), .B(n8), .Y(n1) );
  OR2X2 U3 ( .A(n7), .B(n8), .Y(n2) );
  NAND2X1 U4 ( .A(cmd[1]), .B(n324), .Y(n3) );
  INVX2 U5 ( .A(n217), .Y(n277) );
  INVX2 U6 ( .A(n1), .Y(n4) );
  INVX2 U7 ( .A(n82), .Y(n326) );
  INVX2 U8 ( .A(n18), .Y(n19) );
  INVX2 U12 ( .A(n22), .Y(n23) );
  INVX2 U13 ( .A(n26), .Y(n27) );
  INVX2 U14 ( .A(n33), .Y(n34) );
  INVX2 U15 ( .A(n2), .Y(n5) );
  INVX2 U16 ( .A(n188), .Y(n322) );
  INVX2 U17 ( .A(n83), .Y(n321) );
  INVX2 U18 ( .A(n20), .Y(n21) );
  INVX2 U19 ( .A(n24), .Y(n25) );
  INVX2 U20 ( .A(n10), .Y(n11) );
  INVX2 U21 ( .A(b[2]), .Y(n10) );
  INVX2 U22 ( .A(n12), .Y(n13) );
  INVX2 U23 ( .A(b[3]), .Y(n12) );
  INVX2 U24 ( .A(n16), .Y(n17) );
  INVX2 U25 ( .A(a[1]), .Y(n16) );
  INVX2 U26 ( .A(n8), .Y(n9) );
  INVX2 U27 ( .A(b[1]), .Y(n8) );
  INVX2 U28 ( .A(a[2]), .Y(n18) );
  INVX2 U29 ( .A(a[3]), .Y(n20) );
  INVX2 U30 ( .A(n6), .Y(n7) );
  INVX2 U31 ( .A(b[0]), .Y(n6) );
  INVX2 U32 ( .A(n14), .Y(n15) );
  INVX2 U33 ( .A(b[4]), .Y(n14) );
  INVX2 U34 ( .A(a[4]), .Y(n22) );
  INVX2 U35 ( .A(a[5]), .Y(n24) );
  INVX2 U36 ( .A(a[6]), .Y(n26) );
  INVX2 U37 ( .A(n28), .Y(n32) );
  INVX2 U38 ( .A(a[7]), .Y(n28) );
  INVX2 U39 ( .A(a[15]), .Y(n33) );
  INVX2 U40 ( .A(n186), .Y(n323) );
  INVX2 U41 ( .A(n192), .Y(n327) );
  INVX2 U42 ( .A(n193), .Y(n328) );
  INVX2 U43 ( .A(n187), .Y(n325) );
  NAND2X1 U44 ( .A(n7), .B(n9), .Y(n216) );
  NAND2X1 U45 ( .A(n6), .B(n8), .Y(n217) );
  AOI22X1 U46 ( .A(n275), .B(n339), .C(n277), .D(n342), .Y(n36) );
  NAND2X1 U47 ( .A(n6), .B(n9), .Y(n214) );
  NAND2X1 U48 ( .A(n7), .B(n8), .Y(n215) );
  AOI22X1 U49 ( .A(n278), .B(n287), .C(n276), .D(n341), .Y(n35) );
  AND2X1 U50 ( .A(n36), .B(n35), .Y(n260) );
  NAND3X1 U51 ( .A(n13), .B(n14), .C(n10), .Y(n243) );
  NOR2X1 U52 ( .A(n10), .B(n12), .Y(n240) );
  AND2X1 U53 ( .A(n240), .B(n14), .Y(n213) );
  AOI22X1 U183 ( .A(n275), .B(n33), .C(n277), .D(n289), .Y(n38) );
  AOI22X1 U190 ( .A(n278), .B(n293), .C(n276), .D(n336), .Y(n37) );
  NAND2X1 U191 ( .A(n38), .B(n37), .Y(n229) );
  OAI22X1 U192 ( .A(n17), .B(n215), .C(n19), .D(n214), .Y(n40) );
  OAI22X1 U193 ( .A(a[0]), .B(n217), .C(n21), .D(n216), .Y(n39) );
  NAND3X1 U194 ( .A(n12), .B(n14), .C(n10), .Y(n255) );
  OAI21X1 U195 ( .A(n40), .B(n39), .C(n280), .Y(n41) );
  AOI21X1 U196 ( .A(n213), .B(n229), .C(n284), .Y(n42) );
  OAI21X1 U197 ( .A(n260), .B(n243), .C(n42), .Y(n54) );
  OAI22X1 U198 ( .A(n216), .B(n32), .C(n217), .D(a[4]), .Y(n44) );
  OAI22X1 U199 ( .A(n214), .B(a[6]), .C(n215), .D(n25), .Y(n43) );
  NOR2X1 U200 ( .A(n44), .B(n43), .Y(n231) );
  NAND3X1 U201 ( .A(n12), .B(n14), .C(n11), .Y(n259) );
  OR2X1 U202 ( .A(b[6]), .B(b[5]), .Y(n45) );
  NOR2X1 U203 ( .A(b[15]), .B(n45), .Y(n52) );
  OR2X1 U204 ( .A(b[9]), .B(b[8]), .Y(n46) );
  NOR2X1 U205 ( .A(b[7]), .B(n46), .Y(n51) );
  NOR2X1 U206 ( .A(b[11]), .B(b[10]), .Y(n49) );
  OR2X1 U207 ( .A(b[14]), .B(b[13]), .Y(n47) );
  NOR2X1 U208 ( .A(b[12]), .B(n47), .Y(n48) );
  AND2X1 U209 ( .A(n49), .B(n48), .Y(n50) );
  NAND3X1 U210 ( .A(n52), .B(n51), .C(n50), .Y(n258) );
  NOR2X1 U211 ( .A(n14), .B(n34), .Y(n266) );
  NOR2X1 U212 ( .A(n258), .B(n266), .Y(n254) );
  OAI21X1 U213 ( .A(n231), .B(n259), .C(n254), .Y(n53) );
  NOR2X1 U214 ( .A(n54), .B(n53), .Y(N129) );
  MUX2X1 U215 ( .B(n33), .A(n293), .S(n277), .Y(n201) );
  NAND3X1 U216 ( .A(n282), .B(n279), .C(n201), .Y(n58) );
  NAND2X1 U217 ( .A(n34), .B(n14), .Y(n228) );
  NAND2X1 U218 ( .A(n297), .B(n282), .Y(n69) );
  NAND2X1 U219 ( .A(n298), .B(n13), .Y(n265) );
  AOI22X1 U220 ( .A(n275), .B(n336), .C(n277), .D(n287), .Y(n56) );
  AOI22X1 U221 ( .A(n278), .B(n289), .C(n276), .D(n339), .Y(n55) );
  NAND2X1 U222 ( .A(n56), .B(n55), .Y(n244) );
  NOR2X1 U223 ( .A(n258), .B(n255), .Y(n261) );
  OAI21X1 U224 ( .A(n10), .B(n8), .C(n34), .Y(n202) );
  NAND3X1 U225 ( .A(n15), .B(n12), .C(n282), .Y(n70) );
  AOI22X1 U226 ( .A(n292), .B(n261), .C(n300), .D(n283), .Y(n57) );
  NAND3X1 U227 ( .A(n58), .B(n265), .C(n57), .Y(N139) );
  AOI22X1 U228 ( .A(n275), .B(n293), .C(n277), .D(n339), .Y(n60) );
  AOI22X1 U229 ( .A(n278), .B(n336), .C(n276), .D(n289), .Y(n59) );
  NAND2X1 U230 ( .A(n60), .B(n59), .Y(n224) );
  OAI21X1 U231 ( .A(n10), .B(n6), .C(n300), .Y(n212) );
  AOI22X1 U232 ( .A(n294), .B(n261), .C(n301), .D(n283), .Y(n62) );
  OAI21X1 U233 ( .A(n10), .B(n69), .C(n265), .Y(n61) );
  NAND2X1 U234 ( .A(n62), .B(n299), .Y(N140) );
  NAND2X1 U235 ( .A(n283), .B(n34), .Y(n264) );
  AOI22X1 U236 ( .A(n302), .B(n10), .C(n261), .D(n296), .Y(n63) );
  NAND2X1 U237 ( .A(n63), .B(n299), .Y(N141) );
  NOR2X1 U238 ( .A(n11), .B(n70), .Y(n65) );
  NAND2X1 U239 ( .A(n34), .B(n216), .Y(n267) );
  AOI22X1 U240 ( .A(n276), .B(n293), .C(n277), .D(n336), .Y(n64) );
  OAI21X1 U241 ( .A(n34), .B(n8), .C(n64), .Y(n271) );
  AOI22X1 U242 ( .A(n65), .B(n303), .C(n304), .D(n261), .Y(n66) );
  NAND2X1 U243 ( .A(n66), .B(n299), .Y(N142) );
  NOR2X1 U244 ( .A(n11), .B(n9), .Y(n67) );
  AOI22X1 U245 ( .A(n67), .B(n302), .C(n201), .D(n261), .Y(n68) );
  NAND2X1 U246 ( .A(n68), .B(n299), .Y(N143) );
  NAND3X1 U247 ( .A(n34), .B(n10), .C(n277), .Y(n250) );
  OAI21X1 U248 ( .A(n70), .B(n250), .C(n69), .Y(N144) );
  AOI22X1 U249 ( .A(n275), .B(n289), .C(n277), .D(n341), .Y(n72) );
  AOI22X1 U250 ( .A(n278), .B(n339), .C(n276), .D(n287), .Y(n71) );
  NAND2X1 U251 ( .A(n72), .B(n71), .Y(n270) );
  MUX2X1 U252 ( .B(n304), .A(n303), .S(n15), .Y(n195) );
  OAI22X1 U253 ( .A(n216), .B(a[4]), .C(n217), .D(n17), .Y(n80) );
  OAI22X1 U254 ( .A(n214), .B(n21), .C(n215), .D(a[2]), .Y(n73) );
  OAI21X1 U255 ( .A(n80), .B(n73), .C(n280), .Y(n194) );
  AOI21X1 U256 ( .A(n195), .B(n240), .C(n285), .Y(n196) );
  OAI21X1 U257 ( .A(n290), .B(n243), .C(n196), .Y(n200) );
  OAI22X1 U258 ( .A(n216), .B(a[8]), .C(n217), .D(n25), .Y(n198) );
  OAI22X1 U259 ( .A(n214), .B(n32), .C(n215), .D(a[6]), .Y(n197) );
  NOR2X1 U260 ( .A(n198), .B(n197), .Y(n236) );
  OAI21X1 U261 ( .A(n236), .B(n259), .C(n254), .Y(n199) );
  NOR2X1 U262 ( .A(n200), .B(n199), .Y(N130) );
  NOR2X1 U263 ( .A(n12), .B(n14), .Y(n251) );
  AOI22X1 U264 ( .A(n213), .B(n295), .C(n251), .D(n202), .Y(n206) );
  OAI22X1 U265 ( .A(n21), .B(n215), .C(a[4]), .D(n214), .Y(n204) );
  OAI22X1 U266 ( .A(a[2]), .B(n217), .C(n25), .D(n216), .Y(n203) );
  OAI21X1 U267 ( .A(n204), .B(n203), .C(n280), .Y(n205) );
  NAND2X1 U268 ( .A(n206), .B(n205), .Y(n211) );
  OAI22X1 U269 ( .A(n216), .B(a[9]), .C(n217), .D(n27), .Y(n207) );
  AOI22X1 U270 ( .A(n278), .B(n342), .C(n276), .D(n28), .Y(n208) );
  NAND2X1 U271 ( .A(n286), .B(n208), .Y(n245) );
  AOI22X1 U272 ( .A(n281), .B(n244), .C(n279), .D(n245), .Y(n209) );
  NAND2X1 U273 ( .A(n209), .B(n254), .Y(n210) );
  NOR2X1 U274 ( .A(n211), .B(n210), .Y(N131) );
  AOI22X1 U275 ( .A(n213), .B(n33), .C(n251), .D(n212), .Y(n221) );
  OAI22X1 U276 ( .A(a[4]), .B(n215), .C(n25), .D(n214), .Y(n219) );
  OAI22X1 U277 ( .A(n21), .B(n217), .C(n27), .D(n216), .Y(n218) );
  OAI21X1 U278 ( .A(n219), .B(n218), .C(n280), .Y(n220) );
  NAND2X1 U279 ( .A(n221), .B(n220), .Y(n227) );
  AOI22X1 U280 ( .A(n275), .B(n287), .C(n277), .D(n28), .Y(n223) );
  AOI22X1 U281 ( .A(n278), .B(n341), .C(n276), .D(n342), .Y(n222) );
  NAND2X1 U282 ( .A(n223), .B(n222), .Y(n253) );
  AOI22X1 U283 ( .A(n281), .B(n224), .C(n279), .D(n253), .Y(n225) );
  NAND2X1 U284 ( .A(n225), .B(n254), .Y(n226) );
  NOR2X1 U285 ( .A(n227), .B(n226), .Y(N132) );
  AND2X1 U286 ( .A(n240), .B(n228), .Y(n234) );
  AOI21X1 U287 ( .A(n281), .B(n229), .C(n234), .Y(n230) );
  OAI21X1 U288 ( .A(n260), .B(n259), .C(n230), .Y(n233) );
  OAI21X1 U289 ( .A(n231), .B(n255), .C(n254), .Y(n232) );
  NOR2X1 U290 ( .A(n233), .B(n232), .Y(N133) );
  AOI21X1 U291 ( .A(n251), .B(n267), .C(n234), .Y(n235) );
  OAI21X1 U292 ( .A(n304), .B(n243), .C(n235), .Y(n239) );
  OAI22X1 U293 ( .A(n259), .B(n290), .C(n255), .D(n236), .Y(n237) );
  NAND2X1 U294 ( .A(n291), .B(n254), .Y(n238) );
  NOR2X1 U295 ( .A(n239), .B(n238), .Y(N134) );
  AOI21X1 U296 ( .A(n240), .B(n298), .C(n302), .Y(n249) );
  NOR2X1 U297 ( .A(n11), .B(n14), .Y(n241) );
  NAND3X1 U298 ( .A(n34), .B(n8), .C(n241), .Y(n242) );
  OAI21X1 U299 ( .A(n295), .B(n243), .C(n242), .Y(n247) );
  OAI22X1 U300 ( .A(n255), .B(n245), .C(n259), .D(n244), .Y(n246) );
  OAI21X1 U301 ( .A(n247), .B(n246), .C(n282), .Y(n248) );
  NAND2X1 U302 ( .A(n249), .B(n248), .Y(N135) );
  AOI22X1 U303 ( .A(n13), .B(n33), .C(n251), .D(n250), .Y(n252) );
  OAI21X1 U304 ( .A(n294), .B(n259), .C(n252), .Y(n257) );
  OAI21X1 U305 ( .A(n288), .B(n255), .C(n254), .Y(n256) );
  NOR2X1 U306 ( .A(n257), .B(n256), .Y(N136) );
  NOR2X1 U307 ( .A(n259), .B(n258), .Y(n262) );
  AOI22X1 U308 ( .A(n262), .B(n296), .C(n261), .D(n260), .Y(n263) );
  NAND3X1 U309 ( .A(n265), .B(n264), .C(n263), .Y(N137) );
  NOR2X1 U310 ( .A(n14), .B(n10), .Y(n268) );
  AOI21X1 U311 ( .A(n268), .B(n267), .C(n266), .Y(n269) );
  OAI21X1 U312 ( .A(n12), .B(n297), .C(n269), .Y(n274) );
  AOI22X1 U313 ( .A(n279), .B(n271), .C(n280), .D(n270), .Y(n272) );
  NAND2X1 U314 ( .A(n272), .B(n282), .Y(n273) );
  NOR2X1 U315 ( .A(n274), .B(n273), .Y(N138) );
  INVX2 U316 ( .A(n216), .Y(n275) );
  INVX2 U317 ( .A(n215), .Y(n276) );
  INVX2 U318 ( .A(n214), .Y(n278) );
  INVX2 U319 ( .A(n259), .Y(n279) );
  INVX2 U320 ( .A(n255), .Y(n280) );
  INVX2 U321 ( .A(n243), .Y(n281) );
  INVX2 U322 ( .A(n258), .Y(n282) );
  INVX2 U323 ( .A(n70), .Y(n283) );
  INVX2 U324 ( .A(n41), .Y(n284) );
  INVX2 U325 ( .A(n194), .Y(n285) );
  INVX2 U326 ( .A(n207), .Y(n286) );
  INVX2 U327 ( .A(a[10]), .Y(n287) );
  INVX2 U328 ( .A(n253), .Y(n288) );
  INVX2 U329 ( .A(a[12]), .Y(n289) );
  INVX2 U330 ( .A(n270), .Y(n290) );
  INVX2 U331 ( .A(n237), .Y(n291) );
  INVX2 U332 ( .A(n244), .Y(n292) );
  INVX2 U333 ( .A(a[14]), .Y(n293) );
  INVX2 U334 ( .A(n224), .Y(n294) );
  INVX2 U335 ( .A(n201), .Y(n295) );
  INVX2 U336 ( .A(n229), .Y(n296) );
  INVX2 U337 ( .A(n228), .Y(n297) );
  INVX2 U338 ( .A(n69), .Y(n298) );
  INVX2 U339 ( .A(n61), .Y(n299) );
  INVX2 U340 ( .A(n202), .Y(n300) );
  INVX2 U341 ( .A(n212), .Y(n301) );
  INVX2 U342 ( .A(n264), .Y(n302) );
  INVX2 U343 ( .A(n267), .Y(n303) );
  INVX2 U344 ( .A(n271), .Y(n304) );
  OR2X2 U345 ( .A(b[12]), .B(b[11]), .Y(n357) );
  OR2X2 U346 ( .A(b[15]), .B(b[14]), .Y(n358) );
  OR2X2 U347 ( .A(b[6]), .B(b[5]), .Y(n359) );
  OR2X2 U348 ( .A(b[9]), .B(b[8]), .Y(n360) );
  OR2X2 U349 ( .A(n431), .B(n348), .Y(n380) );
  INVX2 U350 ( .A(n143), .Y(n305) );
  INVX2 U351 ( .A(n150), .Y(n306) );
  INVX2 U352 ( .A(n157), .Y(n307) );
  INVX2 U353 ( .A(n164), .Y(n308) );
  INVX2 U354 ( .A(n171), .Y(n309) );
  INVX2 U355 ( .A(n178), .Y(n310) );
  INVX2 U356 ( .A(n77), .Y(n311) );
  INVX2 U357 ( .A(n87), .Y(n312) );
  INVX2 U358 ( .A(n94), .Y(n313) );
  INVX2 U359 ( .A(n101), .Y(n314) );
  INVX2 U360 ( .A(n108), .Y(n315) );
  INVX2 U361 ( .A(n115), .Y(n316) );
  INVX2 U362 ( .A(n122), .Y(n317) );
  INVX2 U363 ( .A(n129), .Y(n318) );
  INVX2 U364 ( .A(n136), .Y(n319) );
  INVX2 U365 ( .A(n185), .Y(n320) );
  INVX2 U366 ( .A(cmd[2]), .Y(n324) );
  INVX2 U367 ( .A(cmd[1]), .Y(n329) );
  INVX2 U368 ( .A(cmd[0]), .Y(n330) );
  INVX2 U369 ( .A(n428), .Y(n331) );
  INVX2 U370 ( .A(n419), .Y(n332) );
  INVX2 U371 ( .A(n416), .Y(n333) );
  INVX2 U372 ( .A(n424), .Y(n334) );
  INVX2 U373 ( .A(n391), .Y(n335) );
  INVX2 U374 ( .A(a[13]), .Y(n336) );
  INVX2 U375 ( .A(n432), .Y(n337) );
  INVX2 U376 ( .A(n429), .Y(n338) );
  INVX2 U377 ( .A(a[11]), .Y(n339) );
  INVX2 U378 ( .A(n427), .Y(n340) );
  INVX2 U379 ( .A(a[9]), .Y(n341) );
  INVX2 U380 ( .A(a[8]), .Y(n342) );
  INVX2 U381 ( .A(n354), .Y(n343) );
  INVX2 U382 ( .A(a[0]), .Y(n344) );
  INVX2 U383 ( .A(n412), .Y(n345) );
  INVX2 U384 ( .A(n430), .Y(n346) );
  INVX2 U385 ( .A(n404), .Y(n347) );
  INVX2 U386 ( .A(n423), .Y(n348) );
  INVX2 U387 ( .A(n401), .Y(n349) );
  NOR2X1 U388 ( .A(n7), .B(n9), .Y(n423) );
  AOI22X1 U389 ( .A(n4), .B(n339), .C(n423), .D(n342), .Y(n351) );
  NOR2X1 U390 ( .A(n6), .B(n9), .Y(n401) );
  AOI22X1 U391 ( .A(n401), .B(n341), .C(n5), .D(n287), .Y(n350) );
  NAND2X1 U392 ( .A(n351), .B(n350), .Y(n429) );
  NAND2X1 U393 ( .A(n13), .B(n10), .Y(n413) );
  NOR2X1 U394 ( .A(n12), .B(n10), .Y(n394) );
  AOI22X1 U395 ( .A(n4), .B(n33), .C(n423), .D(n289), .Y(n353) );
  AOI22X1 U396 ( .A(n401), .B(n336), .C(n5), .D(n293), .Y(n352) );
  NAND2X1 U397 ( .A(n353), .B(n352), .Y(n428) );
  NOR2X1 U398 ( .A(n13), .B(n10), .Y(n404) );
  OAI22X1 U399 ( .A(n1), .B(n32), .C(n348), .D(n23), .Y(n354) );
  AOI22X1 U400 ( .A(n401), .B(n24), .C(n5), .D(n26), .Y(n355) );
  NAND2X1 U401 ( .A(n343), .B(n355), .Y(n415) );
  AOI22X1 U402 ( .A(n394), .B(n428), .C(n404), .D(n415), .Y(n356) );
  OAI21X1 U403 ( .A(n338), .B(n413), .C(n356), .Y(n370) );
  NOR2X1 U404 ( .A(b[10]), .B(n357), .Y(n365) );
  NOR2X1 U405 ( .A(b[13]), .B(n358), .Y(n364) );
  NOR2X1 U406 ( .A(n15), .B(n359), .Y(n362) );
  NOR2X1 U407 ( .A(b[7]), .B(n360), .Y(n361) );
  AND2X1 U408 ( .A(n362), .B(n361), .Y(n363) );
  NAND3X1 U409 ( .A(n365), .B(n364), .C(n363), .Y(n412) );
  OAI22X1 U410 ( .A(a[2]), .B(n2), .C(n17), .D(n349), .Y(n367) );
  OAI22X1 U411 ( .A(a[0]), .B(n348), .C(n21), .D(n1), .Y(n366) );
  NOR2X1 U412 ( .A(n13), .B(n11), .Y(n405) );
  OAI21X1 U413 ( .A(n367), .B(n366), .C(n405), .Y(n368) );
  NAND2X1 U414 ( .A(n345), .B(n368), .Y(n369) );
  NOR2X1 U415 ( .A(n370), .B(n369), .Y(N145) );
  NOR2X1 U416 ( .A(n412), .B(n13), .Y(n377) );
  NAND2X1 U417 ( .A(n377), .B(n10), .Y(n431) );
  AOI22X1 U418 ( .A(n4), .B(n336), .C(n423), .D(n287), .Y(n372) );
  AOI22X1 U419 ( .A(n401), .B(n339), .C(n5), .D(n289), .Y(n371) );
  NAND2X1 U420 ( .A(n372), .B(n371), .Y(n391) );
  NAND2X1 U421 ( .A(n377), .B(n11), .Y(n430) );
  MUX2X1 U422 ( .B(n33), .A(n293), .S(n6), .Y(n373) );
  NAND2X1 U423 ( .A(n373), .B(n8), .Y(n419) );
  OAI22X1 U424 ( .A(n431), .B(n391), .C(n430), .D(n419), .Y(N155) );
  NAND2X1 U425 ( .A(n34), .B(n423), .Y(n376) );
  AOI22X1 U426 ( .A(n4), .B(n293), .C(n423), .D(n339), .Y(n375) );
  AOI22X1 U427 ( .A(n401), .B(n289), .C(n5), .D(n336), .Y(n374) );
  NAND2X1 U428 ( .A(n375), .B(n374), .Y(n424) );
  MUX2X1 U429 ( .B(n376), .A(n424), .S(n10), .Y(n409) );
  AND2X1 U430 ( .A(n377), .B(n409), .Y(N156) );
  NOR2X1 U431 ( .A(n431), .B(n428), .Y(N157) );
  OAI21X1 U432 ( .A(a[13]), .B(n348), .C(n1), .Y(n379) );
  OAI22X1 U433 ( .A(n34), .B(n8), .C(a[14]), .D(n6), .Y(n378) );
  NOR2X1 U434 ( .A(n379), .B(n378), .Y(n416) );
  NOR2X1 U435 ( .A(n333), .B(n431), .Y(N158) );
  NOR2X1 U436 ( .A(n431), .B(n419), .Y(N159) );
  NOR2X1 U437 ( .A(n33), .B(n380), .Y(N160) );
  AOI22X1 U438 ( .A(n4), .B(n289), .C(n423), .D(n341), .Y(n382) );
  AOI22X1 U439 ( .A(n401), .B(n287), .C(n5), .D(n339), .Y(n381) );
  NAND2X1 U440 ( .A(n382), .B(n381), .Y(n432) );
  AOI22X1 U441 ( .A(n4), .B(n342), .C(n423), .D(n24), .Y(n384) );
  AOI22X1 U442 ( .A(n401), .B(n26), .C(n5), .D(n28), .Y(n383) );
  NAND2X1 U443 ( .A(n384), .B(n383), .Y(n418) );
  AOI22X1 U444 ( .A(n394), .B(n333), .C(n404), .D(n418), .Y(n385) );
  OAI21X1 U445 ( .A(n337), .B(n413), .C(n385), .Y(n390) );
  OAI22X1 U446 ( .A(n21), .B(n2), .C(a[2]), .D(n349), .Y(n387) );
  OAI22X1 U447 ( .A(n17), .B(n348), .C(a[4]), .D(n1), .Y(n386) );
  OAI21X1 U448 ( .A(n387), .B(n386), .C(n405), .Y(n388) );
  NAND2X1 U449 ( .A(n345), .B(n388), .Y(n389) );
  NOR2X1 U450 ( .A(n390), .B(n389), .Y(N146) );
  AOI22X1 U451 ( .A(n4), .B(n341), .C(n423), .D(n26), .Y(n393) );
  AOI22X1 U452 ( .A(n401), .B(n28), .C(n5), .D(n342), .Y(n392) );
  NAND2X1 U453 ( .A(n393), .B(n392), .Y(n421) );
  AOI22X1 U454 ( .A(n394), .B(n419), .C(n404), .D(n421), .Y(n395) );
  OAI21X1 U455 ( .A(n335), .B(n413), .C(n395), .Y(n400) );
  OAI22X1 U456 ( .A(a[4]), .B(n2), .C(n21), .D(n349), .Y(n397) );
  OAI22X1 U457 ( .A(a[2]), .B(n348), .C(n25), .D(n1), .Y(n396) );
  OAI21X1 U458 ( .A(n397), .B(n396), .C(n405), .Y(n398) );
  NAND2X1 U459 ( .A(n345), .B(n398), .Y(n399) );
  NOR2X1 U460 ( .A(n400), .B(n399), .Y(N147) );
  AOI22X1 U461 ( .A(n4), .B(n287), .C(n423), .D(n28), .Y(n403) );
  AOI22X1 U462 ( .A(n401), .B(n342), .C(n5), .D(n341), .Y(n402) );
  NAND2X1 U463 ( .A(n403), .B(n402), .Y(n427) );
  OAI22X1 U464 ( .A(n25), .B(n2), .C(a[4]), .D(n349), .Y(n407) );
  OAI22X1 U465 ( .A(n21), .B(n348), .C(a[6]), .D(n1), .Y(n406) );
  OAI21X1 U466 ( .A(n407), .B(n406), .C(n405), .Y(n408) );
  OAI21X1 U467 ( .A(n340), .B(n347), .C(n408), .Y(n411) );
  OAI21X1 U468 ( .A(n12), .B(n409), .C(n345), .Y(n410) );
  NOR2X1 U469 ( .A(n411), .B(n410), .Y(N148) );
  NOR2X1 U470 ( .A(n413), .B(n412), .Y(n422) );
  AOI22X1 U471 ( .A(n422), .B(n331), .C(n338), .D(n346), .Y(n414) );
  OAI21X1 U472 ( .A(n431), .B(n415), .C(n414), .Y(N149) );
  AOI22X1 U473 ( .A(n422), .B(n416), .C(n337), .D(n346), .Y(n417) );
  OAI21X1 U474 ( .A(n431), .B(n418), .C(n417), .Y(N150) );
  AOI22X1 U475 ( .A(n332), .B(n422), .C(n335), .D(n346), .Y(n420) );
  OAI21X1 U476 ( .A(n431), .B(n421), .C(n420), .Y(N151) );
  AND2X1 U477 ( .A(n423), .B(n422), .Y(n425) );
  AOI22X1 U478 ( .A(n425), .B(a[15]), .C(n334), .D(n346), .Y(n426) );
  OAI21X1 U479 ( .A(n431), .B(n427), .C(n426), .Y(N152) );
  OAI22X1 U480 ( .A(n431), .B(n429), .C(n430), .D(n428), .Y(N153) );
  OAI22X1 U481 ( .A(n432), .B(n431), .C(n333), .D(n430), .Y(N154) );
endmodule


module EX_stage ( clk, rst, pipeline_reg_in, pipeline_reg_out );
  input [57:0] pipeline_reg_in;
  output [38:0] pipeline_reg_out;
  input clk, rst;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, n1;
  wire   [15:0] ex_alu_result;

  DFFPOSX1 pipeline_reg_out_reg_38_ ( .D(N41), .CLK(clk), .Q(
        pipeline_reg_out[38]) );
  DFFPOSX1 pipeline_reg_out_reg_37_ ( .D(N40), .CLK(clk), .Q(
        pipeline_reg_out[37]) );
  DFFPOSX1 pipeline_reg_out_reg_36_ ( .D(N39), .CLK(clk), .Q(
        pipeline_reg_out[36]) );
  DFFPOSX1 pipeline_reg_out_reg_35_ ( .D(N38), .CLK(clk), .Q(
        pipeline_reg_out[35]) );
  DFFPOSX1 pipeline_reg_out_reg_34_ ( .D(N37), .CLK(clk), .Q(
        pipeline_reg_out[34]) );
  DFFPOSX1 pipeline_reg_out_reg_33_ ( .D(N36), .CLK(clk), .Q(
        pipeline_reg_out[33]) );
  DFFPOSX1 pipeline_reg_out_reg_32_ ( .D(N35), .CLK(clk), .Q(
        pipeline_reg_out[32]) );
  DFFPOSX1 pipeline_reg_out_reg_31_ ( .D(N34), .CLK(clk), .Q(
        pipeline_reg_out[31]) );
  DFFPOSX1 pipeline_reg_out_reg_30_ ( .D(N33), .CLK(clk), .Q(
        pipeline_reg_out[30]) );
  DFFPOSX1 pipeline_reg_out_reg_29_ ( .D(N32), .CLK(clk), .Q(
        pipeline_reg_out[29]) );
  DFFPOSX1 pipeline_reg_out_reg_28_ ( .D(N31), .CLK(clk), .Q(
        pipeline_reg_out[28]) );
  DFFPOSX1 pipeline_reg_out_reg_27_ ( .D(N30), .CLK(clk), .Q(
        pipeline_reg_out[27]) );
  DFFPOSX1 pipeline_reg_out_reg_26_ ( .D(N29), .CLK(clk), .Q(
        pipeline_reg_out[26]) );
  DFFPOSX1 pipeline_reg_out_reg_25_ ( .D(N28), .CLK(clk), .Q(
        pipeline_reg_out[25]) );
  DFFPOSX1 pipeline_reg_out_reg_24_ ( .D(N27), .CLK(clk), .Q(
        pipeline_reg_out[24]) );
  DFFPOSX1 pipeline_reg_out_reg_23_ ( .D(N26), .CLK(clk), .Q(
        pipeline_reg_out[23]) );
  DFFPOSX1 pipeline_reg_out_reg_22_ ( .D(N25), .CLK(clk), .Q(
        pipeline_reg_out[22]) );
  DFFPOSX1 pipeline_reg_out_reg_21_ ( .D(N24), .CLK(clk), .Q(
        pipeline_reg_out[21]) );
  DFFPOSX1 pipeline_reg_out_reg_20_ ( .D(N23), .CLK(clk), .Q(
        pipeline_reg_out[20]) );
  DFFPOSX1 pipeline_reg_out_reg_19_ ( .D(N22), .CLK(clk), .Q(
        pipeline_reg_out[19]) );
  DFFPOSX1 pipeline_reg_out_reg_18_ ( .D(N21), .CLK(clk), .Q(
        pipeline_reg_out[18]) );
  DFFPOSX1 pipeline_reg_out_reg_17_ ( .D(N20), .CLK(clk), .Q(
        pipeline_reg_out[17]) );
  DFFPOSX1 pipeline_reg_out_reg_16_ ( .D(N19), .CLK(clk), .Q(
        pipeline_reg_out[16]) );
  DFFPOSX1 pipeline_reg_out_reg_15_ ( .D(N18), .CLK(clk), .Q(
        pipeline_reg_out[15]) );
  DFFPOSX1 pipeline_reg_out_reg_14_ ( .D(N17), .CLK(clk), .Q(
        pipeline_reg_out[14]) );
  DFFPOSX1 pipeline_reg_out_reg_13_ ( .D(N16), .CLK(clk), .Q(
        pipeline_reg_out[13]) );
  DFFPOSX1 pipeline_reg_out_reg_12_ ( .D(N15), .CLK(clk), .Q(
        pipeline_reg_out[12]) );
  DFFPOSX1 pipeline_reg_out_reg_11_ ( .D(N14), .CLK(clk), .Q(
        pipeline_reg_out[11]) );
  DFFPOSX1 pipeline_reg_out_reg_10_ ( .D(N13), .CLK(clk), .Q(
        pipeline_reg_out[10]) );
  DFFPOSX1 pipeline_reg_out_reg_9_ ( .D(N12), .CLK(clk), .Q(
        pipeline_reg_out[9]) );
  DFFPOSX1 pipeline_reg_out_reg_8_ ( .D(N11), .CLK(clk), .Q(
        pipeline_reg_out[8]) );
  DFFPOSX1 pipeline_reg_out_reg_7_ ( .D(N10), .CLK(clk), .Q(
        pipeline_reg_out[7]) );
  DFFPOSX1 pipeline_reg_out_reg_6_ ( .D(N9), .CLK(clk), .Q(pipeline_reg_out[6]) );
  DFFPOSX1 pipeline_reg_out_reg_5_ ( .D(N8), .CLK(clk), .Q(pipeline_reg_out[5]) );
  DFFPOSX1 pipeline_reg_out_reg_4_ ( .D(N7), .CLK(clk), .Q(pipeline_reg_out[4]) );
  DFFPOSX1 pipeline_reg_out_reg_3_ ( .D(N6), .CLK(clk), .Q(pipeline_reg_out[3]) );
  DFFPOSX1 pipeline_reg_out_reg_2_ ( .D(N5), .CLK(clk), .Q(pipeline_reg_out[2]) );
  DFFPOSX1 pipeline_reg_out_reg_1_ ( .D(N4), .CLK(clk), .Q(pipeline_reg_out[1]) );
  DFFPOSX1 pipeline_reg_out_reg_0_ ( .D(N3), .CLK(clk), .Q(pipeline_reg_out[0]) );
  AND2X1 U4 ( .A(pipeline_reg_in[6]), .B(n1), .Y(N9) );
  AND2X1 U5 ( .A(pipeline_reg_in[5]), .B(n1), .Y(N8) );
  AND2X1 U6 ( .A(pipeline_reg_in[4]), .B(n1), .Y(N7) );
  AND2X1 U7 ( .A(pipeline_reg_in[3]), .B(n1), .Y(N6) );
  AND2X1 U8 ( .A(pipeline_reg_in[2]), .B(n1), .Y(N5) );
  AND2X1 U9 ( .A(pipeline_reg_in[57]), .B(n1), .Y(N41) );
  AND2X1 U10 ( .A(ex_alu_result[15]), .B(n1), .Y(N40) );
  AND2X1 U11 ( .A(pipeline_reg_in[1]), .B(n1), .Y(N4) );
  AND2X1 U12 ( .A(ex_alu_result[14]), .B(n1), .Y(N39) );
  AND2X1 U13 ( .A(ex_alu_result[13]), .B(n1), .Y(N38) );
  AND2X1 U14 ( .A(ex_alu_result[12]), .B(n1), .Y(N37) );
  AND2X1 U15 ( .A(ex_alu_result[11]), .B(n1), .Y(N36) );
  AND2X1 U16 ( .A(ex_alu_result[10]), .B(n1), .Y(N35) );
  AND2X1 U17 ( .A(ex_alu_result[9]), .B(n1), .Y(N34) );
  AND2X1 U18 ( .A(ex_alu_result[8]), .B(n1), .Y(N33) );
  AND2X1 U19 ( .A(ex_alu_result[7]), .B(n1), .Y(N32) );
  AND2X1 U20 ( .A(ex_alu_result[6]), .B(n1), .Y(N31) );
  AND2X1 U21 ( .A(ex_alu_result[5]), .B(n1), .Y(N30) );
  AND2X1 U22 ( .A(pipeline_reg_in[0]), .B(n1), .Y(N3) );
  AND2X1 U23 ( .A(ex_alu_result[4]), .B(n1), .Y(N29) );
  AND2X1 U24 ( .A(ex_alu_result[3]), .B(n1), .Y(N28) );
  AND2X1 U25 ( .A(ex_alu_result[2]), .B(n1), .Y(N27) );
  AND2X1 U26 ( .A(ex_alu_result[1]), .B(n1), .Y(N26) );
  AND2X1 U27 ( .A(ex_alu_result[0]), .B(n1), .Y(N25) );
  AND2X1 U28 ( .A(pipeline_reg_in[21]), .B(n1), .Y(N24) );
  AND2X1 U29 ( .A(pipeline_reg_in[20]), .B(n1), .Y(N23) );
  AND2X1 U30 ( .A(pipeline_reg_in[19]), .B(n1), .Y(N22) );
  AND2X1 U31 ( .A(pipeline_reg_in[18]), .B(n1), .Y(N21) );
  AND2X1 U32 ( .A(pipeline_reg_in[17]), .B(n1), .Y(N20) );
  AND2X1 U33 ( .A(pipeline_reg_in[16]), .B(n1), .Y(N19) );
  AND2X1 U34 ( .A(pipeline_reg_in[15]), .B(n1), .Y(N18) );
  AND2X1 U35 ( .A(pipeline_reg_in[14]), .B(n1), .Y(N17) );
  AND2X1 U36 ( .A(pipeline_reg_in[13]), .B(n1), .Y(N16) );
  AND2X1 U37 ( .A(pipeline_reg_in[12]), .B(n1), .Y(N15) );
  AND2X1 U38 ( .A(pipeline_reg_in[11]), .B(n1), .Y(N14) );
  AND2X1 U39 ( .A(pipeline_reg_in[10]), .B(n1), .Y(N13) );
  AND2X1 U40 ( .A(pipeline_reg_in[9]), .B(n1), .Y(N12) );
  AND2X1 U41 ( .A(pipeline_reg_in[8]), .B(n1), .Y(N11) );
  AND2X1 U42 ( .A(pipeline_reg_in[7]), .B(n1), .Y(N10) );
  alu alu_inst ( .a(pipeline_reg_in[53:38]), .b(pipeline_reg_in[37:22]), .cmd(
        pipeline_reg_in[56:54]), .r(ex_alu_result) );
  INVX2 U3 ( .A(rst), .Y(n1) );
endmodule


module data_mem ( clk, mem_access_addr, mem_write_data, mem_write_en, 
        mem_read_data );
  input [15:0] mem_access_addr;
  input [15:0] mem_write_data;
  output [15:0] mem_read_data;
  input clk, mem_write_en;
  wire   n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n55, n73, n91, n109, n127, n145, n163, n181, n199, n217,
         n235, n253, n271, n289, n307, n328, n345, n362, n379, n396, n413,
         n430, n447, n464, n481, n498, n515, n532, n549, n566, n583, n602,
         n619, n636, n653, n670, n687, n704, n721, n738, n755, n772, n789,
         n806, n823, n840, n857, n876, n893, n910, n927, n944, n961, n978,
         n995, n1012, n1029, n1046, n1063, n1080, n1097, n1114, n1131, n1150,
         n1167, n1184, n1201, n1218, n1235, n1252, n1269, n1286, n1303, n1320,
         n1337, n1354, n1371, n1388, n1405, n1424, n1441, n1458, n1475, n1492,
         n1509, n1526, n1543, n1560, n1577, n1594, n1611, n1628, n1645, n1662,
         n1679, n1697, n1714, n1731, n1748, n1765, n1782, n1799, n1816, n1833,
         n1850, n1867, n1884, n1901, n1918, n1935, n1952, n1970, n1987, n2004,
         n2021, n2038, n2055, n2072, n2089, n2106, n2123, n2140, n2157, n2174,
         n2191, n2208, n2225, n2243, n2260, n2277, n2294, n2311, n2328, n2345,
         n2362, n2379, n2396, n2413, n2430, n2447, n2464, n2481, n2498, n2517,
         n2534, n2551, n2568, n2585, n2602, n2619, n2636, n2653, n2670, n2687,
         n2704, n2721, n2738, n2755, n2772, n2790, n2807, n2824, n2841, n2858,
         n2875, n2892, n2909, n2926, n2943, n2960, n2977, n2994, n3011, n3028,
         n3045, n3063, n3080, n3097, n3114, n3131, n3148, n3165, n3182, n3199,
         n3216, n3233, n3250, n3267, n3284, n3301, n3318, n3336, n3353, n3370,
         n3387, n3404, n3421, n3438, n3455, n3472, n3489, n3506, n3523, n3540,
         n3557, n3574, n3591, n3610, n3627, n3644, n3661, n3678, n3695, n3712,
         n3729, n3746, n3763, n3780, n3797, n3814, n3831, n3848, n3865, n3883,
         n3900, n3917, n3934, n3951, n3968, n3985, n4002, n4019, n4036, n4053,
         n4070, n4087, n4104, n4121, n4138, n4156, n4175, n4193, n4211, n4229,
         n4247, n4264, n4281, n4298, n4316, n4333, n4350, n4367, n4385, n4402,
         n4419, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071;
  wire   [4095:0] ram;

  DFFPOSX1 ram_reg_255__15_ ( .D(n8532), .CLK(clk), .Q(ram[4095]) );
  DFFPOSX1 ram_reg_255__14_ ( .D(n8531), .CLK(clk), .Q(ram[4094]) );
  DFFPOSX1 ram_reg_255__13_ ( .D(n8530), .CLK(clk), .Q(ram[4093]) );
  DFFPOSX1 ram_reg_255__12_ ( .D(n8529), .CLK(clk), .Q(ram[4092]) );
  DFFPOSX1 ram_reg_255__11_ ( .D(n8528), .CLK(clk), .Q(ram[4091]) );
  DFFPOSX1 ram_reg_255__10_ ( .D(n8527), .CLK(clk), .Q(ram[4090]) );
  DFFPOSX1 ram_reg_255__9_ ( .D(n8526), .CLK(clk), .Q(ram[4089]) );
  DFFPOSX1 ram_reg_255__8_ ( .D(n8525), .CLK(clk), .Q(ram[4088]) );
  DFFPOSX1 ram_reg_255__7_ ( .D(n8524), .CLK(clk), .Q(ram[4087]) );
  DFFPOSX1 ram_reg_255__6_ ( .D(n8523), .CLK(clk), .Q(ram[4086]) );
  DFFPOSX1 ram_reg_255__5_ ( .D(n8522), .CLK(clk), .Q(ram[4085]) );
  DFFPOSX1 ram_reg_255__4_ ( .D(n8521), .CLK(clk), .Q(ram[4084]) );
  DFFPOSX1 ram_reg_255__3_ ( .D(n8520), .CLK(clk), .Q(ram[4083]) );
  DFFPOSX1 ram_reg_255__2_ ( .D(n8519), .CLK(clk), .Q(ram[4082]) );
  DFFPOSX1 ram_reg_255__1_ ( .D(n8518), .CLK(clk), .Q(ram[4081]) );
  DFFPOSX1 ram_reg_255__0_ ( .D(n8517), .CLK(clk), .Q(ram[4080]) );
  DFFPOSX1 ram_reg_254__15_ ( .D(n8516), .CLK(clk), .Q(ram[4079]) );
  DFFPOSX1 ram_reg_254__14_ ( .D(n8515), .CLK(clk), .Q(ram[4078]) );
  DFFPOSX1 ram_reg_254__13_ ( .D(n8514), .CLK(clk), .Q(ram[4077]) );
  DFFPOSX1 ram_reg_254__12_ ( .D(n8513), .CLK(clk), .Q(ram[4076]) );
  DFFPOSX1 ram_reg_254__11_ ( .D(n8512), .CLK(clk), .Q(ram[4075]) );
  DFFPOSX1 ram_reg_254__10_ ( .D(n8511), .CLK(clk), .Q(ram[4074]) );
  DFFPOSX1 ram_reg_254__9_ ( .D(n8510), .CLK(clk), .Q(ram[4073]) );
  DFFPOSX1 ram_reg_254__8_ ( .D(n8509), .CLK(clk), .Q(ram[4072]) );
  DFFPOSX1 ram_reg_254__7_ ( .D(n8508), .CLK(clk), .Q(ram[4071]) );
  DFFPOSX1 ram_reg_254__6_ ( .D(n8507), .CLK(clk), .Q(ram[4070]) );
  DFFPOSX1 ram_reg_254__5_ ( .D(n8506), .CLK(clk), .Q(ram[4069]) );
  DFFPOSX1 ram_reg_254__4_ ( .D(n8505), .CLK(clk), .Q(ram[4068]) );
  DFFPOSX1 ram_reg_254__3_ ( .D(n8504), .CLK(clk), .Q(ram[4067]) );
  DFFPOSX1 ram_reg_254__2_ ( .D(n8503), .CLK(clk), .Q(ram[4066]) );
  DFFPOSX1 ram_reg_254__1_ ( .D(n8502), .CLK(clk), .Q(ram[4065]) );
  DFFPOSX1 ram_reg_254__0_ ( .D(n8501), .CLK(clk), .Q(ram[4064]) );
  DFFPOSX1 ram_reg_253__15_ ( .D(n8500), .CLK(clk), .Q(ram[4063]) );
  DFFPOSX1 ram_reg_253__14_ ( .D(n8499), .CLK(clk), .Q(ram[4062]) );
  DFFPOSX1 ram_reg_253__13_ ( .D(n8498), .CLK(clk), .Q(ram[4061]) );
  DFFPOSX1 ram_reg_253__12_ ( .D(n8497), .CLK(clk), .Q(ram[4060]) );
  DFFPOSX1 ram_reg_253__11_ ( .D(n8496), .CLK(clk), .Q(ram[4059]) );
  DFFPOSX1 ram_reg_253__10_ ( .D(n8495), .CLK(clk), .Q(ram[4058]) );
  DFFPOSX1 ram_reg_253__9_ ( .D(n8494), .CLK(clk), .Q(ram[4057]) );
  DFFPOSX1 ram_reg_253__8_ ( .D(n8493), .CLK(clk), .Q(ram[4056]) );
  DFFPOSX1 ram_reg_253__7_ ( .D(n8492), .CLK(clk), .Q(ram[4055]) );
  DFFPOSX1 ram_reg_253__6_ ( .D(n8491), .CLK(clk), .Q(ram[4054]) );
  DFFPOSX1 ram_reg_253__5_ ( .D(n8490), .CLK(clk), .Q(ram[4053]) );
  DFFPOSX1 ram_reg_253__4_ ( .D(n8489), .CLK(clk), .Q(ram[4052]) );
  DFFPOSX1 ram_reg_253__3_ ( .D(n8488), .CLK(clk), .Q(ram[4051]) );
  DFFPOSX1 ram_reg_253__2_ ( .D(n8487), .CLK(clk), .Q(ram[4050]) );
  DFFPOSX1 ram_reg_253__1_ ( .D(n8486), .CLK(clk), .Q(ram[4049]) );
  DFFPOSX1 ram_reg_253__0_ ( .D(n8485), .CLK(clk), .Q(ram[4048]) );
  DFFPOSX1 ram_reg_252__15_ ( .D(n8484), .CLK(clk), .Q(ram[4047]) );
  DFFPOSX1 ram_reg_252__14_ ( .D(n8483), .CLK(clk), .Q(ram[4046]) );
  DFFPOSX1 ram_reg_252__13_ ( .D(n8482), .CLK(clk), .Q(ram[4045]) );
  DFFPOSX1 ram_reg_252__12_ ( .D(n8481), .CLK(clk), .Q(ram[4044]) );
  DFFPOSX1 ram_reg_252__11_ ( .D(n8480), .CLK(clk), .Q(ram[4043]) );
  DFFPOSX1 ram_reg_252__10_ ( .D(n8479), .CLK(clk), .Q(ram[4042]) );
  DFFPOSX1 ram_reg_252__9_ ( .D(n8478), .CLK(clk), .Q(ram[4041]) );
  DFFPOSX1 ram_reg_252__8_ ( .D(n8477), .CLK(clk), .Q(ram[4040]) );
  DFFPOSX1 ram_reg_252__7_ ( .D(n8476), .CLK(clk), .Q(ram[4039]) );
  DFFPOSX1 ram_reg_252__6_ ( .D(n8475), .CLK(clk), .Q(ram[4038]) );
  DFFPOSX1 ram_reg_252__5_ ( .D(n8474), .CLK(clk), .Q(ram[4037]) );
  DFFPOSX1 ram_reg_252__4_ ( .D(n8473), .CLK(clk), .Q(ram[4036]) );
  DFFPOSX1 ram_reg_252__3_ ( .D(n8472), .CLK(clk), .Q(ram[4035]) );
  DFFPOSX1 ram_reg_252__2_ ( .D(n8471), .CLK(clk), .Q(ram[4034]) );
  DFFPOSX1 ram_reg_252__1_ ( .D(n8470), .CLK(clk), .Q(ram[4033]) );
  DFFPOSX1 ram_reg_252__0_ ( .D(n8469), .CLK(clk), .Q(ram[4032]) );
  DFFPOSX1 ram_reg_251__15_ ( .D(n8468), .CLK(clk), .Q(ram[4031]) );
  DFFPOSX1 ram_reg_251__14_ ( .D(n8467), .CLK(clk), .Q(ram[4030]) );
  DFFPOSX1 ram_reg_251__13_ ( .D(n8466), .CLK(clk), .Q(ram[4029]) );
  DFFPOSX1 ram_reg_251__12_ ( .D(n8465), .CLK(clk), .Q(ram[4028]) );
  DFFPOSX1 ram_reg_251__11_ ( .D(n8464), .CLK(clk), .Q(ram[4027]) );
  DFFPOSX1 ram_reg_251__10_ ( .D(n8463), .CLK(clk), .Q(ram[4026]) );
  DFFPOSX1 ram_reg_251__9_ ( .D(n8462), .CLK(clk), .Q(ram[4025]) );
  DFFPOSX1 ram_reg_251__8_ ( .D(n8461), .CLK(clk), .Q(ram[4024]) );
  DFFPOSX1 ram_reg_251__7_ ( .D(n8460), .CLK(clk), .Q(ram[4023]) );
  DFFPOSX1 ram_reg_251__6_ ( .D(n8459), .CLK(clk), .Q(ram[4022]) );
  DFFPOSX1 ram_reg_251__5_ ( .D(n8458), .CLK(clk), .Q(ram[4021]) );
  DFFPOSX1 ram_reg_251__4_ ( .D(n8457), .CLK(clk), .Q(ram[4020]) );
  DFFPOSX1 ram_reg_251__3_ ( .D(n8456), .CLK(clk), .Q(ram[4019]) );
  DFFPOSX1 ram_reg_251__2_ ( .D(n8455), .CLK(clk), .Q(ram[4018]) );
  DFFPOSX1 ram_reg_251__1_ ( .D(n8454), .CLK(clk), .Q(ram[4017]) );
  DFFPOSX1 ram_reg_251__0_ ( .D(n8453), .CLK(clk), .Q(ram[4016]) );
  DFFPOSX1 ram_reg_250__15_ ( .D(n8452), .CLK(clk), .Q(ram[4015]) );
  DFFPOSX1 ram_reg_250__14_ ( .D(n8451), .CLK(clk), .Q(ram[4014]) );
  DFFPOSX1 ram_reg_250__13_ ( .D(n8450), .CLK(clk), .Q(ram[4013]) );
  DFFPOSX1 ram_reg_250__12_ ( .D(n8449), .CLK(clk), .Q(ram[4012]) );
  DFFPOSX1 ram_reg_250__11_ ( .D(n8448), .CLK(clk), .Q(ram[4011]) );
  DFFPOSX1 ram_reg_250__10_ ( .D(n8447), .CLK(clk), .Q(ram[4010]) );
  DFFPOSX1 ram_reg_250__9_ ( .D(n8446), .CLK(clk), .Q(ram[4009]) );
  DFFPOSX1 ram_reg_250__8_ ( .D(n8445), .CLK(clk), .Q(ram[4008]) );
  DFFPOSX1 ram_reg_250__7_ ( .D(n8444), .CLK(clk), .Q(ram[4007]) );
  DFFPOSX1 ram_reg_250__6_ ( .D(n8443), .CLK(clk), .Q(ram[4006]) );
  DFFPOSX1 ram_reg_250__5_ ( .D(n8442), .CLK(clk), .Q(ram[4005]) );
  DFFPOSX1 ram_reg_250__4_ ( .D(n8441), .CLK(clk), .Q(ram[4004]) );
  DFFPOSX1 ram_reg_250__3_ ( .D(n8440), .CLK(clk), .Q(ram[4003]) );
  DFFPOSX1 ram_reg_250__2_ ( .D(n8439), .CLK(clk), .Q(ram[4002]) );
  DFFPOSX1 ram_reg_250__1_ ( .D(n8438), .CLK(clk), .Q(ram[4001]) );
  DFFPOSX1 ram_reg_250__0_ ( .D(n8437), .CLK(clk), .Q(ram[4000]) );
  DFFPOSX1 ram_reg_249__15_ ( .D(n8436), .CLK(clk), .Q(ram[3999]) );
  DFFPOSX1 ram_reg_249__14_ ( .D(n8435), .CLK(clk), .Q(ram[3998]) );
  DFFPOSX1 ram_reg_249__13_ ( .D(n8434), .CLK(clk), .Q(ram[3997]) );
  DFFPOSX1 ram_reg_249__12_ ( .D(n8433), .CLK(clk), .Q(ram[3996]) );
  DFFPOSX1 ram_reg_249__11_ ( .D(n8432), .CLK(clk), .Q(ram[3995]) );
  DFFPOSX1 ram_reg_249__10_ ( .D(n8431), .CLK(clk), .Q(ram[3994]) );
  DFFPOSX1 ram_reg_249__9_ ( .D(n8430), .CLK(clk), .Q(ram[3993]) );
  DFFPOSX1 ram_reg_249__8_ ( .D(n8429), .CLK(clk), .Q(ram[3992]) );
  DFFPOSX1 ram_reg_249__7_ ( .D(n8428), .CLK(clk), .Q(ram[3991]) );
  DFFPOSX1 ram_reg_249__6_ ( .D(n8427), .CLK(clk), .Q(ram[3990]) );
  DFFPOSX1 ram_reg_249__5_ ( .D(n8426), .CLK(clk), .Q(ram[3989]) );
  DFFPOSX1 ram_reg_249__4_ ( .D(n8425), .CLK(clk), .Q(ram[3988]) );
  DFFPOSX1 ram_reg_249__3_ ( .D(n8424), .CLK(clk), .Q(ram[3987]) );
  DFFPOSX1 ram_reg_249__2_ ( .D(n8423), .CLK(clk), .Q(ram[3986]) );
  DFFPOSX1 ram_reg_249__1_ ( .D(n8422), .CLK(clk), .Q(ram[3985]) );
  DFFPOSX1 ram_reg_249__0_ ( .D(n8421), .CLK(clk), .Q(ram[3984]) );
  DFFPOSX1 ram_reg_248__15_ ( .D(n8420), .CLK(clk), .Q(ram[3983]) );
  DFFPOSX1 ram_reg_248__14_ ( .D(n8419), .CLK(clk), .Q(ram[3982]) );
  DFFPOSX1 ram_reg_248__13_ ( .D(n8418), .CLK(clk), .Q(ram[3981]) );
  DFFPOSX1 ram_reg_248__12_ ( .D(n8417), .CLK(clk), .Q(ram[3980]) );
  DFFPOSX1 ram_reg_248__11_ ( .D(n8416), .CLK(clk), .Q(ram[3979]) );
  DFFPOSX1 ram_reg_248__10_ ( .D(n8415), .CLK(clk), .Q(ram[3978]) );
  DFFPOSX1 ram_reg_248__9_ ( .D(n8414), .CLK(clk), .Q(ram[3977]) );
  DFFPOSX1 ram_reg_248__8_ ( .D(n8413), .CLK(clk), .Q(ram[3976]) );
  DFFPOSX1 ram_reg_248__7_ ( .D(n8412), .CLK(clk), .Q(ram[3975]) );
  DFFPOSX1 ram_reg_248__6_ ( .D(n8411), .CLK(clk), .Q(ram[3974]) );
  DFFPOSX1 ram_reg_248__5_ ( .D(n8410), .CLK(clk), .Q(ram[3973]) );
  DFFPOSX1 ram_reg_248__4_ ( .D(n8409), .CLK(clk), .Q(ram[3972]) );
  DFFPOSX1 ram_reg_248__3_ ( .D(n8408), .CLK(clk), .Q(ram[3971]) );
  DFFPOSX1 ram_reg_248__2_ ( .D(n8407), .CLK(clk), .Q(ram[3970]) );
  DFFPOSX1 ram_reg_248__1_ ( .D(n8406), .CLK(clk), .Q(ram[3969]) );
  DFFPOSX1 ram_reg_248__0_ ( .D(n8405), .CLK(clk), .Q(ram[3968]) );
  DFFPOSX1 ram_reg_247__15_ ( .D(n8404), .CLK(clk), .Q(ram[3967]) );
  DFFPOSX1 ram_reg_247__14_ ( .D(n8403), .CLK(clk), .Q(ram[3966]) );
  DFFPOSX1 ram_reg_247__13_ ( .D(n8402), .CLK(clk), .Q(ram[3965]) );
  DFFPOSX1 ram_reg_247__12_ ( .D(n8401), .CLK(clk), .Q(ram[3964]) );
  DFFPOSX1 ram_reg_247__11_ ( .D(n8400), .CLK(clk), .Q(ram[3963]) );
  DFFPOSX1 ram_reg_247__10_ ( .D(n8399), .CLK(clk), .Q(ram[3962]) );
  DFFPOSX1 ram_reg_247__9_ ( .D(n8398), .CLK(clk), .Q(ram[3961]) );
  DFFPOSX1 ram_reg_247__8_ ( .D(n8397), .CLK(clk), .Q(ram[3960]) );
  DFFPOSX1 ram_reg_247__7_ ( .D(n8396), .CLK(clk), .Q(ram[3959]) );
  DFFPOSX1 ram_reg_247__6_ ( .D(n8395), .CLK(clk), .Q(ram[3958]) );
  DFFPOSX1 ram_reg_247__5_ ( .D(n8394), .CLK(clk), .Q(ram[3957]) );
  DFFPOSX1 ram_reg_247__4_ ( .D(n8393), .CLK(clk), .Q(ram[3956]) );
  DFFPOSX1 ram_reg_247__3_ ( .D(n8392), .CLK(clk), .Q(ram[3955]) );
  DFFPOSX1 ram_reg_247__2_ ( .D(n8391), .CLK(clk), .Q(ram[3954]) );
  DFFPOSX1 ram_reg_247__1_ ( .D(n8390), .CLK(clk), .Q(ram[3953]) );
  DFFPOSX1 ram_reg_247__0_ ( .D(n8389), .CLK(clk), .Q(ram[3952]) );
  DFFPOSX1 ram_reg_246__15_ ( .D(n8388), .CLK(clk), .Q(ram[3951]) );
  DFFPOSX1 ram_reg_246__14_ ( .D(n8387), .CLK(clk), .Q(ram[3950]) );
  DFFPOSX1 ram_reg_246__13_ ( .D(n8386), .CLK(clk), .Q(ram[3949]) );
  DFFPOSX1 ram_reg_246__12_ ( .D(n8385), .CLK(clk), .Q(ram[3948]) );
  DFFPOSX1 ram_reg_246__11_ ( .D(n8384), .CLK(clk), .Q(ram[3947]) );
  DFFPOSX1 ram_reg_246__10_ ( .D(n8383), .CLK(clk), .Q(ram[3946]) );
  DFFPOSX1 ram_reg_246__9_ ( .D(n8382), .CLK(clk), .Q(ram[3945]) );
  DFFPOSX1 ram_reg_246__8_ ( .D(n8381), .CLK(clk), .Q(ram[3944]) );
  DFFPOSX1 ram_reg_246__7_ ( .D(n8380), .CLK(clk), .Q(ram[3943]) );
  DFFPOSX1 ram_reg_246__6_ ( .D(n8379), .CLK(clk), .Q(ram[3942]) );
  DFFPOSX1 ram_reg_246__5_ ( .D(n8378), .CLK(clk), .Q(ram[3941]) );
  DFFPOSX1 ram_reg_246__4_ ( .D(n8377), .CLK(clk), .Q(ram[3940]) );
  DFFPOSX1 ram_reg_246__3_ ( .D(n8376), .CLK(clk), .Q(ram[3939]) );
  DFFPOSX1 ram_reg_246__2_ ( .D(n8375), .CLK(clk), .Q(ram[3938]) );
  DFFPOSX1 ram_reg_246__1_ ( .D(n8374), .CLK(clk), .Q(ram[3937]) );
  DFFPOSX1 ram_reg_246__0_ ( .D(n8373), .CLK(clk), .Q(ram[3936]) );
  DFFPOSX1 ram_reg_245__15_ ( .D(n8372), .CLK(clk), .Q(ram[3935]) );
  DFFPOSX1 ram_reg_245__14_ ( .D(n8371), .CLK(clk), .Q(ram[3934]) );
  DFFPOSX1 ram_reg_245__13_ ( .D(n8370), .CLK(clk), .Q(ram[3933]) );
  DFFPOSX1 ram_reg_245__12_ ( .D(n8369), .CLK(clk), .Q(ram[3932]) );
  DFFPOSX1 ram_reg_245__11_ ( .D(n8368), .CLK(clk), .Q(ram[3931]) );
  DFFPOSX1 ram_reg_245__10_ ( .D(n8367), .CLK(clk), .Q(ram[3930]) );
  DFFPOSX1 ram_reg_245__9_ ( .D(n8366), .CLK(clk), .Q(ram[3929]) );
  DFFPOSX1 ram_reg_245__8_ ( .D(n8365), .CLK(clk), .Q(ram[3928]) );
  DFFPOSX1 ram_reg_245__7_ ( .D(n8364), .CLK(clk), .Q(ram[3927]) );
  DFFPOSX1 ram_reg_245__6_ ( .D(n8363), .CLK(clk), .Q(ram[3926]) );
  DFFPOSX1 ram_reg_245__5_ ( .D(n8362), .CLK(clk), .Q(ram[3925]) );
  DFFPOSX1 ram_reg_245__4_ ( .D(n8361), .CLK(clk), .Q(ram[3924]) );
  DFFPOSX1 ram_reg_245__3_ ( .D(n8360), .CLK(clk), .Q(ram[3923]) );
  DFFPOSX1 ram_reg_245__2_ ( .D(n8359), .CLK(clk), .Q(ram[3922]) );
  DFFPOSX1 ram_reg_245__1_ ( .D(n8358), .CLK(clk), .Q(ram[3921]) );
  DFFPOSX1 ram_reg_245__0_ ( .D(n8357), .CLK(clk), .Q(ram[3920]) );
  DFFPOSX1 ram_reg_244__15_ ( .D(n8356), .CLK(clk), .Q(ram[3919]) );
  DFFPOSX1 ram_reg_244__14_ ( .D(n8355), .CLK(clk), .Q(ram[3918]) );
  DFFPOSX1 ram_reg_244__13_ ( .D(n8354), .CLK(clk), .Q(ram[3917]) );
  DFFPOSX1 ram_reg_244__12_ ( .D(n8353), .CLK(clk), .Q(ram[3916]) );
  DFFPOSX1 ram_reg_244__11_ ( .D(n8352), .CLK(clk), .Q(ram[3915]) );
  DFFPOSX1 ram_reg_244__10_ ( .D(n8351), .CLK(clk), .Q(ram[3914]) );
  DFFPOSX1 ram_reg_244__9_ ( .D(n8350), .CLK(clk), .Q(ram[3913]) );
  DFFPOSX1 ram_reg_244__8_ ( .D(n8349), .CLK(clk), .Q(ram[3912]) );
  DFFPOSX1 ram_reg_244__7_ ( .D(n8348), .CLK(clk), .Q(ram[3911]) );
  DFFPOSX1 ram_reg_244__6_ ( .D(n8347), .CLK(clk), .Q(ram[3910]) );
  DFFPOSX1 ram_reg_244__5_ ( .D(n8346), .CLK(clk), .Q(ram[3909]) );
  DFFPOSX1 ram_reg_244__4_ ( .D(n8345), .CLK(clk), .Q(ram[3908]) );
  DFFPOSX1 ram_reg_244__3_ ( .D(n8344), .CLK(clk), .Q(ram[3907]) );
  DFFPOSX1 ram_reg_244__2_ ( .D(n8343), .CLK(clk), .Q(ram[3906]) );
  DFFPOSX1 ram_reg_244__1_ ( .D(n8342), .CLK(clk), .Q(ram[3905]) );
  DFFPOSX1 ram_reg_244__0_ ( .D(n8341), .CLK(clk), .Q(ram[3904]) );
  DFFPOSX1 ram_reg_243__15_ ( .D(n8340), .CLK(clk), .Q(ram[3903]) );
  DFFPOSX1 ram_reg_243__14_ ( .D(n8339), .CLK(clk), .Q(ram[3902]) );
  DFFPOSX1 ram_reg_243__13_ ( .D(n8338), .CLK(clk), .Q(ram[3901]) );
  DFFPOSX1 ram_reg_243__12_ ( .D(n8337), .CLK(clk), .Q(ram[3900]) );
  DFFPOSX1 ram_reg_243__11_ ( .D(n8336), .CLK(clk), .Q(ram[3899]) );
  DFFPOSX1 ram_reg_243__10_ ( .D(n8335), .CLK(clk), .Q(ram[3898]) );
  DFFPOSX1 ram_reg_243__9_ ( .D(n8334), .CLK(clk), .Q(ram[3897]) );
  DFFPOSX1 ram_reg_243__8_ ( .D(n8333), .CLK(clk), .Q(ram[3896]) );
  DFFPOSX1 ram_reg_243__7_ ( .D(n8332), .CLK(clk), .Q(ram[3895]) );
  DFFPOSX1 ram_reg_243__6_ ( .D(n8331), .CLK(clk), .Q(ram[3894]) );
  DFFPOSX1 ram_reg_243__5_ ( .D(n8330), .CLK(clk), .Q(ram[3893]) );
  DFFPOSX1 ram_reg_243__4_ ( .D(n8329), .CLK(clk), .Q(ram[3892]) );
  DFFPOSX1 ram_reg_243__3_ ( .D(n8328), .CLK(clk), .Q(ram[3891]) );
  DFFPOSX1 ram_reg_243__2_ ( .D(n8327), .CLK(clk), .Q(ram[3890]) );
  DFFPOSX1 ram_reg_243__1_ ( .D(n8326), .CLK(clk), .Q(ram[3889]) );
  DFFPOSX1 ram_reg_243__0_ ( .D(n8325), .CLK(clk), .Q(ram[3888]) );
  DFFPOSX1 ram_reg_242__15_ ( .D(n8324), .CLK(clk), .Q(ram[3887]) );
  DFFPOSX1 ram_reg_242__14_ ( .D(n8323), .CLK(clk), .Q(ram[3886]) );
  DFFPOSX1 ram_reg_242__13_ ( .D(n8322), .CLK(clk), .Q(ram[3885]) );
  DFFPOSX1 ram_reg_242__12_ ( .D(n8321), .CLK(clk), .Q(ram[3884]) );
  DFFPOSX1 ram_reg_242__11_ ( .D(n8320), .CLK(clk), .Q(ram[3883]) );
  DFFPOSX1 ram_reg_242__10_ ( .D(n8319), .CLK(clk), .Q(ram[3882]) );
  DFFPOSX1 ram_reg_242__9_ ( .D(n8318), .CLK(clk), .Q(ram[3881]) );
  DFFPOSX1 ram_reg_242__8_ ( .D(n8317), .CLK(clk), .Q(ram[3880]) );
  DFFPOSX1 ram_reg_242__7_ ( .D(n8316), .CLK(clk), .Q(ram[3879]) );
  DFFPOSX1 ram_reg_242__6_ ( .D(n8315), .CLK(clk), .Q(ram[3878]) );
  DFFPOSX1 ram_reg_242__5_ ( .D(n8314), .CLK(clk), .Q(ram[3877]) );
  DFFPOSX1 ram_reg_242__4_ ( .D(n8313), .CLK(clk), .Q(ram[3876]) );
  DFFPOSX1 ram_reg_242__3_ ( .D(n8312), .CLK(clk), .Q(ram[3875]) );
  DFFPOSX1 ram_reg_242__2_ ( .D(n8311), .CLK(clk), .Q(ram[3874]) );
  DFFPOSX1 ram_reg_242__1_ ( .D(n8310), .CLK(clk), .Q(ram[3873]) );
  DFFPOSX1 ram_reg_242__0_ ( .D(n8309), .CLK(clk), .Q(ram[3872]) );
  DFFPOSX1 ram_reg_241__15_ ( .D(n8308), .CLK(clk), .Q(ram[3871]) );
  DFFPOSX1 ram_reg_241__14_ ( .D(n8307), .CLK(clk), .Q(ram[3870]) );
  DFFPOSX1 ram_reg_241__13_ ( .D(n8306), .CLK(clk), .Q(ram[3869]) );
  DFFPOSX1 ram_reg_241__12_ ( .D(n8305), .CLK(clk), .Q(ram[3868]) );
  DFFPOSX1 ram_reg_241__11_ ( .D(n8304), .CLK(clk), .Q(ram[3867]) );
  DFFPOSX1 ram_reg_241__10_ ( .D(n8303), .CLK(clk), .Q(ram[3866]) );
  DFFPOSX1 ram_reg_241__9_ ( .D(n8302), .CLK(clk), .Q(ram[3865]) );
  DFFPOSX1 ram_reg_241__8_ ( .D(n8301), .CLK(clk), .Q(ram[3864]) );
  DFFPOSX1 ram_reg_241__7_ ( .D(n8300), .CLK(clk), .Q(ram[3863]) );
  DFFPOSX1 ram_reg_241__6_ ( .D(n8299), .CLK(clk), .Q(ram[3862]) );
  DFFPOSX1 ram_reg_241__5_ ( .D(n8298), .CLK(clk), .Q(ram[3861]) );
  DFFPOSX1 ram_reg_241__4_ ( .D(n8297), .CLK(clk), .Q(ram[3860]) );
  DFFPOSX1 ram_reg_241__3_ ( .D(n8296), .CLK(clk), .Q(ram[3859]) );
  DFFPOSX1 ram_reg_241__2_ ( .D(n8295), .CLK(clk), .Q(ram[3858]) );
  DFFPOSX1 ram_reg_241__1_ ( .D(n8294), .CLK(clk), .Q(ram[3857]) );
  DFFPOSX1 ram_reg_241__0_ ( .D(n8293), .CLK(clk), .Q(ram[3856]) );
  DFFPOSX1 ram_reg_240__15_ ( .D(n8292), .CLK(clk), .Q(ram[3855]) );
  DFFPOSX1 ram_reg_240__14_ ( .D(n8291), .CLK(clk), .Q(ram[3854]) );
  DFFPOSX1 ram_reg_240__13_ ( .D(n8290), .CLK(clk), .Q(ram[3853]) );
  DFFPOSX1 ram_reg_240__12_ ( .D(n8289), .CLK(clk), .Q(ram[3852]) );
  DFFPOSX1 ram_reg_240__11_ ( .D(n8288), .CLK(clk), .Q(ram[3851]) );
  DFFPOSX1 ram_reg_240__10_ ( .D(n8287), .CLK(clk), .Q(ram[3850]) );
  DFFPOSX1 ram_reg_240__9_ ( .D(n8286), .CLK(clk), .Q(ram[3849]) );
  DFFPOSX1 ram_reg_240__8_ ( .D(n8285), .CLK(clk), .Q(ram[3848]) );
  DFFPOSX1 ram_reg_240__7_ ( .D(n8284), .CLK(clk), .Q(ram[3847]) );
  DFFPOSX1 ram_reg_240__6_ ( .D(n8283), .CLK(clk), .Q(ram[3846]) );
  DFFPOSX1 ram_reg_240__5_ ( .D(n8282), .CLK(clk), .Q(ram[3845]) );
  DFFPOSX1 ram_reg_240__4_ ( .D(n8281), .CLK(clk), .Q(ram[3844]) );
  DFFPOSX1 ram_reg_240__3_ ( .D(n8280), .CLK(clk), .Q(ram[3843]) );
  DFFPOSX1 ram_reg_240__2_ ( .D(n8279), .CLK(clk), .Q(ram[3842]) );
  DFFPOSX1 ram_reg_240__1_ ( .D(n8278), .CLK(clk), .Q(ram[3841]) );
  DFFPOSX1 ram_reg_240__0_ ( .D(n8277), .CLK(clk), .Q(ram[3840]) );
  DFFPOSX1 ram_reg_239__15_ ( .D(n8276), .CLK(clk), .Q(ram[3839]) );
  DFFPOSX1 ram_reg_239__14_ ( .D(n8275), .CLK(clk), .Q(ram[3838]) );
  DFFPOSX1 ram_reg_239__13_ ( .D(n8274), .CLK(clk), .Q(ram[3837]) );
  DFFPOSX1 ram_reg_239__12_ ( .D(n8273), .CLK(clk), .Q(ram[3836]) );
  DFFPOSX1 ram_reg_239__11_ ( .D(n8272), .CLK(clk), .Q(ram[3835]) );
  DFFPOSX1 ram_reg_239__10_ ( .D(n8271), .CLK(clk), .Q(ram[3834]) );
  DFFPOSX1 ram_reg_239__9_ ( .D(n8270), .CLK(clk), .Q(ram[3833]) );
  DFFPOSX1 ram_reg_239__8_ ( .D(n8269), .CLK(clk), .Q(ram[3832]) );
  DFFPOSX1 ram_reg_239__7_ ( .D(n8268), .CLK(clk), .Q(ram[3831]) );
  DFFPOSX1 ram_reg_239__6_ ( .D(n8267), .CLK(clk), .Q(ram[3830]) );
  DFFPOSX1 ram_reg_239__5_ ( .D(n8266), .CLK(clk), .Q(ram[3829]) );
  DFFPOSX1 ram_reg_239__4_ ( .D(n8265), .CLK(clk), .Q(ram[3828]) );
  DFFPOSX1 ram_reg_239__3_ ( .D(n8264), .CLK(clk), .Q(ram[3827]) );
  DFFPOSX1 ram_reg_239__2_ ( .D(n8263), .CLK(clk), .Q(ram[3826]) );
  DFFPOSX1 ram_reg_239__1_ ( .D(n8262), .CLK(clk), .Q(ram[3825]) );
  DFFPOSX1 ram_reg_239__0_ ( .D(n8261), .CLK(clk), .Q(ram[3824]) );
  DFFPOSX1 ram_reg_238__15_ ( .D(n8260), .CLK(clk), .Q(ram[3823]) );
  DFFPOSX1 ram_reg_238__14_ ( .D(n8259), .CLK(clk), .Q(ram[3822]) );
  DFFPOSX1 ram_reg_238__13_ ( .D(n8258), .CLK(clk), .Q(ram[3821]) );
  DFFPOSX1 ram_reg_238__12_ ( .D(n8257), .CLK(clk), .Q(ram[3820]) );
  DFFPOSX1 ram_reg_238__11_ ( .D(n8256), .CLK(clk), .Q(ram[3819]) );
  DFFPOSX1 ram_reg_238__10_ ( .D(n8255), .CLK(clk), .Q(ram[3818]) );
  DFFPOSX1 ram_reg_238__9_ ( .D(n8254), .CLK(clk), .Q(ram[3817]) );
  DFFPOSX1 ram_reg_238__8_ ( .D(n8253), .CLK(clk), .Q(ram[3816]) );
  DFFPOSX1 ram_reg_238__7_ ( .D(n8252), .CLK(clk), .Q(ram[3815]) );
  DFFPOSX1 ram_reg_238__6_ ( .D(n8251), .CLK(clk), .Q(ram[3814]) );
  DFFPOSX1 ram_reg_238__5_ ( .D(n8250), .CLK(clk), .Q(ram[3813]) );
  DFFPOSX1 ram_reg_238__4_ ( .D(n8249), .CLK(clk), .Q(ram[3812]) );
  DFFPOSX1 ram_reg_238__3_ ( .D(n8248), .CLK(clk), .Q(ram[3811]) );
  DFFPOSX1 ram_reg_238__2_ ( .D(n8247), .CLK(clk), .Q(ram[3810]) );
  DFFPOSX1 ram_reg_238__1_ ( .D(n8246), .CLK(clk), .Q(ram[3809]) );
  DFFPOSX1 ram_reg_238__0_ ( .D(n8245), .CLK(clk), .Q(ram[3808]) );
  DFFPOSX1 ram_reg_237__15_ ( .D(n8244), .CLK(clk), .Q(ram[3807]) );
  DFFPOSX1 ram_reg_237__14_ ( .D(n8243), .CLK(clk), .Q(ram[3806]) );
  DFFPOSX1 ram_reg_237__13_ ( .D(n8242), .CLK(clk), .Q(ram[3805]) );
  DFFPOSX1 ram_reg_237__12_ ( .D(n8241), .CLK(clk), .Q(ram[3804]) );
  DFFPOSX1 ram_reg_237__11_ ( .D(n8240), .CLK(clk), .Q(ram[3803]) );
  DFFPOSX1 ram_reg_237__10_ ( .D(n8239), .CLK(clk), .Q(ram[3802]) );
  DFFPOSX1 ram_reg_237__9_ ( .D(n8238), .CLK(clk), .Q(ram[3801]) );
  DFFPOSX1 ram_reg_237__8_ ( .D(n8237), .CLK(clk), .Q(ram[3800]) );
  DFFPOSX1 ram_reg_237__7_ ( .D(n8236), .CLK(clk), .Q(ram[3799]) );
  DFFPOSX1 ram_reg_237__6_ ( .D(n8235), .CLK(clk), .Q(ram[3798]) );
  DFFPOSX1 ram_reg_237__5_ ( .D(n8234), .CLK(clk), .Q(ram[3797]) );
  DFFPOSX1 ram_reg_237__4_ ( .D(n8233), .CLK(clk), .Q(ram[3796]) );
  DFFPOSX1 ram_reg_237__3_ ( .D(n8232), .CLK(clk), .Q(ram[3795]) );
  DFFPOSX1 ram_reg_237__2_ ( .D(n8231), .CLK(clk), .Q(ram[3794]) );
  DFFPOSX1 ram_reg_237__1_ ( .D(n8230), .CLK(clk), .Q(ram[3793]) );
  DFFPOSX1 ram_reg_237__0_ ( .D(n8229), .CLK(clk), .Q(ram[3792]) );
  DFFPOSX1 ram_reg_236__15_ ( .D(n8228), .CLK(clk), .Q(ram[3791]) );
  DFFPOSX1 ram_reg_236__14_ ( .D(n8227), .CLK(clk), .Q(ram[3790]) );
  DFFPOSX1 ram_reg_236__13_ ( .D(n8226), .CLK(clk), .Q(ram[3789]) );
  DFFPOSX1 ram_reg_236__12_ ( .D(n8225), .CLK(clk), .Q(ram[3788]) );
  DFFPOSX1 ram_reg_236__11_ ( .D(n8224), .CLK(clk), .Q(ram[3787]) );
  DFFPOSX1 ram_reg_236__10_ ( .D(n8223), .CLK(clk), .Q(ram[3786]) );
  DFFPOSX1 ram_reg_236__9_ ( .D(n8222), .CLK(clk), .Q(ram[3785]) );
  DFFPOSX1 ram_reg_236__8_ ( .D(n8221), .CLK(clk), .Q(ram[3784]) );
  DFFPOSX1 ram_reg_236__7_ ( .D(n8220), .CLK(clk), .Q(ram[3783]) );
  DFFPOSX1 ram_reg_236__6_ ( .D(n8219), .CLK(clk), .Q(ram[3782]) );
  DFFPOSX1 ram_reg_236__5_ ( .D(n8218), .CLK(clk), .Q(ram[3781]) );
  DFFPOSX1 ram_reg_236__4_ ( .D(n8217), .CLK(clk), .Q(ram[3780]) );
  DFFPOSX1 ram_reg_236__3_ ( .D(n8216), .CLK(clk), .Q(ram[3779]) );
  DFFPOSX1 ram_reg_236__2_ ( .D(n8215), .CLK(clk), .Q(ram[3778]) );
  DFFPOSX1 ram_reg_236__1_ ( .D(n8214), .CLK(clk), .Q(ram[3777]) );
  DFFPOSX1 ram_reg_236__0_ ( .D(n8213), .CLK(clk), .Q(ram[3776]) );
  DFFPOSX1 ram_reg_235__15_ ( .D(n8212), .CLK(clk), .Q(ram[3775]) );
  DFFPOSX1 ram_reg_235__14_ ( .D(n8211), .CLK(clk), .Q(ram[3774]) );
  DFFPOSX1 ram_reg_235__13_ ( .D(n8210), .CLK(clk), .Q(ram[3773]) );
  DFFPOSX1 ram_reg_235__12_ ( .D(n8209), .CLK(clk), .Q(ram[3772]) );
  DFFPOSX1 ram_reg_235__11_ ( .D(n8208), .CLK(clk), .Q(ram[3771]) );
  DFFPOSX1 ram_reg_235__10_ ( .D(n8207), .CLK(clk), .Q(ram[3770]) );
  DFFPOSX1 ram_reg_235__9_ ( .D(n8206), .CLK(clk), .Q(ram[3769]) );
  DFFPOSX1 ram_reg_235__8_ ( .D(n8205), .CLK(clk), .Q(ram[3768]) );
  DFFPOSX1 ram_reg_235__7_ ( .D(n8204), .CLK(clk), .Q(ram[3767]) );
  DFFPOSX1 ram_reg_235__6_ ( .D(n8203), .CLK(clk), .Q(ram[3766]) );
  DFFPOSX1 ram_reg_235__5_ ( .D(n8202), .CLK(clk), .Q(ram[3765]) );
  DFFPOSX1 ram_reg_235__4_ ( .D(n8201), .CLK(clk), .Q(ram[3764]) );
  DFFPOSX1 ram_reg_235__3_ ( .D(n8200), .CLK(clk), .Q(ram[3763]) );
  DFFPOSX1 ram_reg_235__2_ ( .D(n8199), .CLK(clk), .Q(ram[3762]) );
  DFFPOSX1 ram_reg_235__1_ ( .D(n8198), .CLK(clk), .Q(ram[3761]) );
  DFFPOSX1 ram_reg_235__0_ ( .D(n8197), .CLK(clk), .Q(ram[3760]) );
  DFFPOSX1 ram_reg_234__15_ ( .D(n8196), .CLK(clk), .Q(ram[3759]) );
  DFFPOSX1 ram_reg_234__14_ ( .D(n8195), .CLK(clk), .Q(ram[3758]) );
  DFFPOSX1 ram_reg_234__13_ ( .D(n8194), .CLK(clk), .Q(ram[3757]) );
  DFFPOSX1 ram_reg_234__12_ ( .D(n8193), .CLK(clk), .Q(ram[3756]) );
  DFFPOSX1 ram_reg_234__11_ ( .D(n8192), .CLK(clk), .Q(ram[3755]) );
  DFFPOSX1 ram_reg_234__10_ ( .D(n8191), .CLK(clk), .Q(ram[3754]) );
  DFFPOSX1 ram_reg_234__9_ ( .D(n8190), .CLK(clk), .Q(ram[3753]) );
  DFFPOSX1 ram_reg_234__8_ ( .D(n8189), .CLK(clk), .Q(ram[3752]) );
  DFFPOSX1 ram_reg_234__7_ ( .D(n8188), .CLK(clk), .Q(ram[3751]) );
  DFFPOSX1 ram_reg_234__6_ ( .D(n8187), .CLK(clk), .Q(ram[3750]) );
  DFFPOSX1 ram_reg_234__5_ ( .D(n8186), .CLK(clk), .Q(ram[3749]) );
  DFFPOSX1 ram_reg_234__4_ ( .D(n8185), .CLK(clk), .Q(ram[3748]) );
  DFFPOSX1 ram_reg_234__3_ ( .D(n8184), .CLK(clk), .Q(ram[3747]) );
  DFFPOSX1 ram_reg_234__2_ ( .D(n8183), .CLK(clk), .Q(ram[3746]) );
  DFFPOSX1 ram_reg_234__1_ ( .D(n8182), .CLK(clk), .Q(ram[3745]) );
  DFFPOSX1 ram_reg_234__0_ ( .D(n8181), .CLK(clk), .Q(ram[3744]) );
  DFFPOSX1 ram_reg_233__15_ ( .D(n8180), .CLK(clk), .Q(ram[3743]) );
  DFFPOSX1 ram_reg_233__14_ ( .D(n8179), .CLK(clk), .Q(ram[3742]) );
  DFFPOSX1 ram_reg_233__13_ ( .D(n8178), .CLK(clk), .Q(ram[3741]) );
  DFFPOSX1 ram_reg_233__12_ ( .D(n8177), .CLK(clk), .Q(ram[3740]) );
  DFFPOSX1 ram_reg_233__11_ ( .D(n8176), .CLK(clk), .Q(ram[3739]) );
  DFFPOSX1 ram_reg_233__10_ ( .D(n8175), .CLK(clk), .Q(ram[3738]) );
  DFFPOSX1 ram_reg_233__9_ ( .D(n8174), .CLK(clk), .Q(ram[3737]) );
  DFFPOSX1 ram_reg_233__8_ ( .D(n8173), .CLK(clk), .Q(ram[3736]) );
  DFFPOSX1 ram_reg_233__7_ ( .D(n8172), .CLK(clk), .Q(ram[3735]) );
  DFFPOSX1 ram_reg_233__6_ ( .D(n8171), .CLK(clk), .Q(ram[3734]) );
  DFFPOSX1 ram_reg_233__5_ ( .D(n8170), .CLK(clk), .Q(ram[3733]) );
  DFFPOSX1 ram_reg_233__4_ ( .D(n8169), .CLK(clk), .Q(ram[3732]) );
  DFFPOSX1 ram_reg_233__3_ ( .D(n8168), .CLK(clk), .Q(ram[3731]) );
  DFFPOSX1 ram_reg_233__2_ ( .D(n8167), .CLK(clk), .Q(ram[3730]) );
  DFFPOSX1 ram_reg_233__1_ ( .D(n8166), .CLK(clk), .Q(ram[3729]) );
  DFFPOSX1 ram_reg_233__0_ ( .D(n8165), .CLK(clk), .Q(ram[3728]) );
  DFFPOSX1 ram_reg_232__15_ ( .D(n8164), .CLK(clk), .Q(ram[3727]) );
  DFFPOSX1 ram_reg_232__14_ ( .D(n8163), .CLK(clk), .Q(ram[3726]) );
  DFFPOSX1 ram_reg_232__13_ ( .D(n8162), .CLK(clk), .Q(ram[3725]) );
  DFFPOSX1 ram_reg_232__12_ ( .D(n8161), .CLK(clk), .Q(ram[3724]) );
  DFFPOSX1 ram_reg_232__11_ ( .D(n8160), .CLK(clk), .Q(ram[3723]) );
  DFFPOSX1 ram_reg_232__10_ ( .D(n8159), .CLK(clk), .Q(ram[3722]) );
  DFFPOSX1 ram_reg_232__9_ ( .D(n8158), .CLK(clk), .Q(ram[3721]) );
  DFFPOSX1 ram_reg_232__8_ ( .D(n8157), .CLK(clk), .Q(ram[3720]) );
  DFFPOSX1 ram_reg_232__7_ ( .D(n8156), .CLK(clk), .Q(ram[3719]) );
  DFFPOSX1 ram_reg_232__6_ ( .D(n8155), .CLK(clk), .Q(ram[3718]) );
  DFFPOSX1 ram_reg_232__5_ ( .D(n8154), .CLK(clk), .Q(ram[3717]) );
  DFFPOSX1 ram_reg_232__4_ ( .D(n8153), .CLK(clk), .Q(ram[3716]) );
  DFFPOSX1 ram_reg_232__3_ ( .D(n8152), .CLK(clk), .Q(ram[3715]) );
  DFFPOSX1 ram_reg_232__2_ ( .D(n8151), .CLK(clk), .Q(ram[3714]) );
  DFFPOSX1 ram_reg_232__1_ ( .D(n8150), .CLK(clk), .Q(ram[3713]) );
  DFFPOSX1 ram_reg_232__0_ ( .D(n8149), .CLK(clk), .Q(ram[3712]) );
  DFFPOSX1 ram_reg_231__15_ ( .D(n8148), .CLK(clk), .Q(ram[3711]) );
  DFFPOSX1 ram_reg_231__14_ ( .D(n8147), .CLK(clk), .Q(ram[3710]) );
  DFFPOSX1 ram_reg_231__13_ ( .D(n8146), .CLK(clk), .Q(ram[3709]) );
  DFFPOSX1 ram_reg_231__12_ ( .D(n8145), .CLK(clk), .Q(ram[3708]) );
  DFFPOSX1 ram_reg_231__11_ ( .D(n8144), .CLK(clk), .Q(ram[3707]) );
  DFFPOSX1 ram_reg_231__10_ ( .D(n8143), .CLK(clk), .Q(ram[3706]) );
  DFFPOSX1 ram_reg_231__9_ ( .D(n8142), .CLK(clk), .Q(ram[3705]) );
  DFFPOSX1 ram_reg_231__8_ ( .D(n8141), .CLK(clk), .Q(ram[3704]) );
  DFFPOSX1 ram_reg_231__7_ ( .D(n8140), .CLK(clk), .Q(ram[3703]) );
  DFFPOSX1 ram_reg_231__6_ ( .D(n8139), .CLK(clk), .Q(ram[3702]) );
  DFFPOSX1 ram_reg_231__5_ ( .D(n8138), .CLK(clk), .Q(ram[3701]) );
  DFFPOSX1 ram_reg_231__4_ ( .D(n8137), .CLK(clk), .Q(ram[3700]) );
  DFFPOSX1 ram_reg_231__3_ ( .D(n8136), .CLK(clk), .Q(ram[3699]) );
  DFFPOSX1 ram_reg_231__2_ ( .D(n8135), .CLK(clk), .Q(ram[3698]) );
  DFFPOSX1 ram_reg_231__1_ ( .D(n8134), .CLK(clk), .Q(ram[3697]) );
  DFFPOSX1 ram_reg_231__0_ ( .D(n8133), .CLK(clk), .Q(ram[3696]) );
  DFFPOSX1 ram_reg_230__15_ ( .D(n8132), .CLK(clk), .Q(ram[3695]) );
  DFFPOSX1 ram_reg_230__14_ ( .D(n8131), .CLK(clk), .Q(ram[3694]) );
  DFFPOSX1 ram_reg_230__13_ ( .D(n8130), .CLK(clk), .Q(ram[3693]) );
  DFFPOSX1 ram_reg_230__12_ ( .D(n8129), .CLK(clk), .Q(ram[3692]) );
  DFFPOSX1 ram_reg_230__11_ ( .D(n8128), .CLK(clk), .Q(ram[3691]) );
  DFFPOSX1 ram_reg_230__10_ ( .D(n8127), .CLK(clk), .Q(ram[3690]) );
  DFFPOSX1 ram_reg_230__9_ ( .D(n8126), .CLK(clk), .Q(ram[3689]) );
  DFFPOSX1 ram_reg_230__8_ ( .D(n8125), .CLK(clk), .Q(ram[3688]) );
  DFFPOSX1 ram_reg_230__7_ ( .D(n8124), .CLK(clk), .Q(ram[3687]) );
  DFFPOSX1 ram_reg_230__6_ ( .D(n8123), .CLK(clk), .Q(ram[3686]) );
  DFFPOSX1 ram_reg_230__5_ ( .D(n8122), .CLK(clk), .Q(ram[3685]) );
  DFFPOSX1 ram_reg_230__4_ ( .D(n8121), .CLK(clk), .Q(ram[3684]) );
  DFFPOSX1 ram_reg_230__3_ ( .D(n8120), .CLK(clk), .Q(ram[3683]) );
  DFFPOSX1 ram_reg_230__2_ ( .D(n8119), .CLK(clk), .Q(ram[3682]) );
  DFFPOSX1 ram_reg_230__1_ ( .D(n8118), .CLK(clk), .Q(ram[3681]) );
  DFFPOSX1 ram_reg_230__0_ ( .D(n8117), .CLK(clk), .Q(ram[3680]) );
  DFFPOSX1 ram_reg_229__15_ ( .D(n8116), .CLK(clk), .Q(ram[3679]) );
  DFFPOSX1 ram_reg_229__14_ ( .D(n8115), .CLK(clk), .Q(ram[3678]) );
  DFFPOSX1 ram_reg_229__13_ ( .D(n8114), .CLK(clk), .Q(ram[3677]) );
  DFFPOSX1 ram_reg_229__12_ ( .D(n8113), .CLK(clk), .Q(ram[3676]) );
  DFFPOSX1 ram_reg_229__11_ ( .D(n8112), .CLK(clk), .Q(ram[3675]) );
  DFFPOSX1 ram_reg_229__10_ ( .D(n8111), .CLK(clk), .Q(ram[3674]) );
  DFFPOSX1 ram_reg_229__9_ ( .D(n8110), .CLK(clk), .Q(ram[3673]) );
  DFFPOSX1 ram_reg_229__8_ ( .D(n8109), .CLK(clk), .Q(ram[3672]) );
  DFFPOSX1 ram_reg_229__7_ ( .D(n8108), .CLK(clk), .Q(ram[3671]) );
  DFFPOSX1 ram_reg_229__6_ ( .D(n8107), .CLK(clk), .Q(ram[3670]) );
  DFFPOSX1 ram_reg_229__5_ ( .D(n8106), .CLK(clk), .Q(ram[3669]) );
  DFFPOSX1 ram_reg_229__4_ ( .D(n8105), .CLK(clk), .Q(ram[3668]) );
  DFFPOSX1 ram_reg_229__3_ ( .D(n8104), .CLK(clk), .Q(ram[3667]) );
  DFFPOSX1 ram_reg_229__2_ ( .D(n8103), .CLK(clk), .Q(ram[3666]) );
  DFFPOSX1 ram_reg_229__1_ ( .D(n8102), .CLK(clk), .Q(ram[3665]) );
  DFFPOSX1 ram_reg_229__0_ ( .D(n8101), .CLK(clk), .Q(ram[3664]) );
  DFFPOSX1 ram_reg_228__15_ ( .D(n8100), .CLK(clk), .Q(ram[3663]) );
  DFFPOSX1 ram_reg_228__14_ ( .D(n8099), .CLK(clk), .Q(ram[3662]) );
  DFFPOSX1 ram_reg_228__13_ ( .D(n8098), .CLK(clk), .Q(ram[3661]) );
  DFFPOSX1 ram_reg_228__12_ ( .D(n8097), .CLK(clk), .Q(ram[3660]) );
  DFFPOSX1 ram_reg_228__11_ ( .D(n8096), .CLK(clk), .Q(ram[3659]) );
  DFFPOSX1 ram_reg_228__10_ ( .D(n8095), .CLK(clk), .Q(ram[3658]) );
  DFFPOSX1 ram_reg_228__9_ ( .D(n8094), .CLK(clk), .Q(ram[3657]) );
  DFFPOSX1 ram_reg_228__8_ ( .D(n8093), .CLK(clk), .Q(ram[3656]) );
  DFFPOSX1 ram_reg_228__7_ ( .D(n8092), .CLK(clk), .Q(ram[3655]) );
  DFFPOSX1 ram_reg_228__6_ ( .D(n8091), .CLK(clk), .Q(ram[3654]) );
  DFFPOSX1 ram_reg_228__5_ ( .D(n8090), .CLK(clk), .Q(ram[3653]) );
  DFFPOSX1 ram_reg_228__4_ ( .D(n8089), .CLK(clk), .Q(ram[3652]) );
  DFFPOSX1 ram_reg_228__3_ ( .D(n8088), .CLK(clk), .Q(ram[3651]) );
  DFFPOSX1 ram_reg_228__2_ ( .D(n8087), .CLK(clk), .Q(ram[3650]) );
  DFFPOSX1 ram_reg_228__1_ ( .D(n8086), .CLK(clk), .Q(ram[3649]) );
  DFFPOSX1 ram_reg_228__0_ ( .D(n8085), .CLK(clk), .Q(ram[3648]) );
  DFFPOSX1 ram_reg_227__15_ ( .D(n8084), .CLK(clk), .Q(ram[3647]) );
  DFFPOSX1 ram_reg_227__14_ ( .D(n8083), .CLK(clk), .Q(ram[3646]) );
  DFFPOSX1 ram_reg_227__13_ ( .D(n8082), .CLK(clk), .Q(ram[3645]) );
  DFFPOSX1 ram_reg_227__12_ ( .D(n8081), .CLK(clk), .Q(ram[3644]) );
  DFFPOSX1 ram_reg_227__11_ ( .D(n8080), .CLK(clk), .Q(ram[3643]) );
  DFFPOSX1 ram_reg_227__10_ ( .D(n8079), .CLK(clk), .Q(ram[3642]) );
  DFFPOSX1 ram_reg_227__9_ ( .D(n8078), .CLK(clk), .Q(ram[3641]) );
  DFFPOSX1 ram_reg_227__8_ ( .D(n8077), .CLK(clk), .Q(ram[3640]) );
  DFFPOSX1 ram_reg_227__7_ ( .D(n8076), .CLK(clk), .Q(ram[3639]) );
  DFFPOSX1 ram_reg_227__6_ ( .D(n8075), .CLK(clk), .Q(ram[3638]) );
  DFFPOSX1 ram_reg_227__5_ ( .D(n8074), .CLK(clk), .Q(ram[3637]) );
  DFFPOSX1 ram_reg_227__4_ ( .D(n8073), .CLK(clk), .Q(ram[3636]) );
  DFFPOSX1 ram_reg_227__3_ ( .D(n8072), .CLK(clk), .Q(ram[3635]) );
  DFFPOSX1 ram_reg_227__2_ ( .D(n8071), .CLK(clk), .Q(ram[3634]) );
  DFFPOSX1 ram_reg_227__1_ ( .D(n8070), .CLK(clk), .Q(ram[3633]) );
  DFFPOSX1 ram_reg_227__0_ ( .D(n8069), .CLK(clk), .Q(ram[3632]) );
  DFFPOSX1 ram_reg_226__15_ ( .D(n8068), .CLK(clk), .Q(ram[3631]) );
  DFFPOSX1 ram_reg_226__14_ ( .D(n8067), .CLK(clk), .Q(ram[3630]) );
  DFFPOSX1 ram_reg_226__13_ ( .D(n8066), .CLK(clk), .Q(ram[3629]) );
  DFFPOSX1 ram_reg_226__12_ ( .D(n8065), .CLK(clk), .Q(ram[3628]) );
  DFFPOSX1 ram_reg_226__11_ ( .D(n8064), .CLK(clk), .Q(ram[3627]) );
  DFFPOSX1 ram_reg_226__10_ ( .D(n8063), .CLK(clk), .Q(ram[3626]) );
  DFFPOSX1 ram_reg_226__9_ ( .D(n8062), .CLK(clk), .Q(ram[3625]) );
  DFFPOSX1 ram_reg_226__8_ ( .D(n8061), .CLK(clk), .Q(ram[3624]) );
  DFFPOSX1 ram_reg_226__7_ ( .D(n8060), .CLK(clk), .Q(ram[3623]) );
  DFFPOSX1 ram_reg_226__6_ ( .D(n8059), .CLK(clk), .Q(ram[3622]) );
  DFFPOSX1 ram_reg_226__5_ ( .D(n8058), .CLK(clk), .Q(ram[3621]) );
  DFFPOSX1 ram_reg_226__4_ ( .D(n8057), .CLK(clk), .Q(ram[3620]) );
  DFFPOSX1 ram_reg_226__3_ ( .D(n8056), .CLK(clk), .Q(ram[3619]) );
  DFFPOSX1 ram_reg_226__2_ ( .D(n8055), .CLK(clk), .Q(ram[3618]) );
  DFFPOSX1 ram_reg_226__1_ ( .D(n8054), .CLK(clk), .Q(ram[3617]) );
  DFFPOSX1 ram_reg_226__0_ ( .D(n8053), .CLK(clk), .Q(ram[3616]) );
  DFFPOSX1 ram_reg_225__15_ ( .D(n8052), .CLK(clk), .Q(ram[3615]) );
  DFFPOSX1 ram_reg_225__14_ ( .D(n8051), .CLK(clk), .Q(ram[3614]) );
  DFFPOSX1 ram_reg_225__13_ ( .D(n8050), .CLK(clk), .Q(ram[3613]) );
  DFFPOSX1 ram_reg_225__12_ ( .D(n8049), .CLK(clk), .Q(ram[3612]) );
  DFFPOSX1 ram_reg_225__11_ ( .D(n8048), .CLK(clk), .Q(ram[3611]) );
  DFFPOSX1 ram_reg_225__10_ ( .D(n8047), .CLK(clk), .Q(ram[3610]) );
  DFFPOSX1 ram_reg_225__9_ ( .D(n8046), .CLK(clk), .Q(ram[3609]) );
  DFFPOSX1 ram_reg_225__8_ ( .D(n8045), .CLK(clk), .Q(ram[3608]) );
  DFFPOSX1 ram_reg_225__7_ ( .D(n8044), .CLK(clk), .Q(ram[3607]) );
  DFFPOSX1 ram_reg_225__6_ ( .D(n8043), .CLK(clk), .Q(ram[3606]) );
  DFFPOSX1 ram_reg_225__5_ ( .D(n8042), .CLK(clk), .Q(ram[3605]) );
  DFFPOSX1 ram_reg_225__4_ ( .D(n8041), .CLK(clk), .Q(ram[3604]) );
  DFFPOSX1 ram_reg_225__3_ ( .D(n8040), .CLK(clk), .Q(ram[3603]) );
  DFFPOSX1 ram_reg_225__2_ ( .D(n8039), .CLK(clk), .Q(ram[3602]) );
  DFFPOSX1 ram_reg_225__1_ ( .D(n8038), .CLK(clk), .Q(ram[3601]) );
  DFFPOSX1 ram_reg_225__0_ ( .D(n8037), .CLK(clk), .Q(ram[3600]) );
  DFFPOSX1 ram_reg_224__15_ ( .D(n8036), .CLK(clk), .Q(ram[3599]) );
  DFFPOSX1 ram_reg_224__14_ ( .D(n8035), .CLK(clk), .Q(ram[3598]) );
  DFFPOSX1 ram_reg_224__13_ ( .D(n8034), .CLK(clk), .Q(ram[3597]) );
  DFFPOSX1 ram_reg_224__12_ ( .D(n8033), .CLK(clk), .Q(ram[3596]) );
  DFFPOSX1 ram_reg_224__11_ ( .D(n8032), .CLK(clk), .Q(ram[3595]) );
  DFFPOSX1 ram_reg_224__10_ ( .D(n8031), .CLK(clk), .Q(ram[3594]) );
  DFFPOSX1 ram_reg_224__9_ ( .D(n8030), .CLK(clk), .Q(ram[3593]) );
  DFFPOSX1 ram_reg_224__8_ ( .D(n8029), .CLK(clk), .Q(ram[3592]) );
  DFFPOSX1 ram_reg_224__7_ ( .D(n8028), .CLK(clk), .Q(ram[3591]) );
  DFFPOSX1 ram_reg_224__6_ ( .D(n8027), .CLK(clk), .Q(ram[3590]) );
  DFFPOSX1 ram_reg_224__5_ ( .D(n8026), .CLK(clk), .Q(ram[3589]) );
  DFFPOSX1 ram_reg_224__4_ ( .D(n8025), .CLK(clk), .Q(ram[3588]) );
  DFFPOSX1 ram_reg_224__3_ ( .D(n8024), .CLK(clk), .Q(ram[3587]) );
  DFFPOSX1 ram_reg_224__2_ ( .D(n8023), .CLK(clk), .Q(ram[3586]) );
  DFFPOSX1 ram_reg_224__1_ ( .D(n8022), .CLK(clk), .Q(ram[3585]) );
  DFFPOSX1 ram_reg_224__0_ ( .D(n8021), .CLK(clk), .Q(ram[3584]) );
  DFFPOSX1 ram_reg_223__15_ ( .D(n8020), .CLK(clk), .Q(ram[3583]) );
  DFFPOSX1 ram_reg_223__14_ ( .D(n8019), .CLK(clk), .Q(ram[3582]) );
  DFFPOSX1 ram_reg_223__13_ ( .D(n8018), .CLK(clk), .Q(ram[3581]) );
  DFFPOSX1 ram_reg_223__12_ ( .D(n8017), .CLK(clk), .Q(ram[3580]) );
  DFFPOSX1 ram_reg_223__11_ ( .D(n8016), .CLK(clk), .Q(ram[3579]) );
  DFFPOSX1 ram_reg_223__10_ ( .D(n8015), .CLK(clk), .Q(ram[3578]) );
  DFFPOSX1 ram_reg_223__9_ ( .D(n8014), .CLK(clk), .Q(ram[3577]) );
  DFFPOSX1 ram_reg_223__8_ ( .D(n8013), .CLK(clk), .Q(ram[3576]) );
  DFFPOSX1 ram_reg_223__7_ ( .D(n8012), .CLK(clk), .Q(ram[3575]) );
  DFFPOSX1 ram_reg_223__6_ ( .D(n8011), .CLK(clk), .Q(ram[3574]) );
  DFFPOSX1 ram_reg_223__5_ ( .D(n8010), .CLK(clk), .Q(ram[3573]) );
  DFFPOSX1 ram_reg_223__4_ ( .D(n8009), .CLK(clk), .Q(ram[3572]) );
  DFFPOSX1 ram_reg_223__3_ ( .D(n8008), .CLK(clk), .Q(ram[3571]) );
  DFFPOSX1 ram_reg_223__2_ ( .D(n8007), .CLK(clk), .Q(ram[3570]) );
  DFFPOSX1 ram_reg_223__1_ ( .D(n8006), .CLK(clk), .Q(ram[3569]) );
  DFFPOSX1 ram_reg_223__0_ ( .D(n8005), .CLK(clk), .Q(ram[3568]) );
  DFFPOSX1 ram_reg_222__15_ ( .D(n8004), .CLK(clk), .Q(ram[3567]) );
  DFFPOSX1 ram_reg_222__14_ ( .D(n8003), .CLK(clk), .Q(ram[3566]) );
  DFFPOSX1 ram_reg_222__13_ ( .D(n8002), .CLK(clk), .Q(ram[3565]) );
  DFFPOSX1 ram_reg_222__12_ ( .D(n8001), .CLK(clk), .Q(ram[3564]) );
  DFFPOSX1 ram_reg_222__11_ ( .D(n8000), .CLK(clk), .Q(ram[3563]) );
  DFFPOSX1 ram_reg_222__10_ ( .D(n7999), .CLK(clk), .Q(ram[3562]) );
  DFFPOSX1 ram_reg_222__9_ ( .D(n7998), .CLK(clk), .Q(ram[3561]) );
  DFFPOSX1 ram_reg_222__8_ ( .D(n7997), .CLK(clk), .Q(ram[3560]) );
  DFFPOSX1 ram_reg_222__7_ ( .D(n7996), .CLK(clk), .Q(ram[3559]) );
  DFFPOSX1 ram_reg_222__6_ ( .D(n7995), .CLK(clk), .Q(ram[3558]) );
  DFFPOSX1 ram_reg_222__5_ ( .D(n7994), .CLK(clk), .Q(ram[3557]) );
  DFFPOSX1 ram_reg_222__4_ ( .D(n7993), .CLK(clk), .Q(ram[3556]) );
  DFFPOSX1 ram_reg_222__3_ ( .D(n7992), .CLK(clk), .Q(ram[3555]) );
  DFFPOSX1 ram_reg_222__2_ ( .D(n7991), .CLK(clk), .Q(ram[3554]) );
  DFFPOSX1 ram_reg_222__1_ ( .D(n7990), .CLK(clk), .Q(ram[3553]) );
  DFFPOSX1 ram_reg_222__0_ ( .D(n7989), .CLK(clk), .Q(ram[3552]) );
  DFFPOSX1 ram_reg_221__15_ ( .D(n7988), .CLK(clk), .Q(ram[3551]) );
  DFFPOSX1 ram_reg_221__14_ ( .D(n7987), .CLK(clk), .Q(ram[3550]) );
  DFFPOSX1 ram_reg_221__13_ ( .D(n7986), .CLK(clk), .Q(ram[3549]) );
  DFFPOSX1 ram_reg_221__12_ ( .D(n7985), .CLK(clk), .Q(ram[3548]) );
  DFFPOSX1 ram_reg_221__11_ ( .D(n7984), .CLK(clk), .Q(ram[3547]) );
  DFFPOSX1 ram_reg_221__10_ ( .D(n7983), .CLK(clk), .Q(ram[3546]) );
  DFFPOSX1 ram_reg_221__9_ ( .D(n7982), .CLK(clk), .Q(ram[3545]) );
  DFFPOSX1 ram_reg_221__8_ ( .D(n7981), .CLK(clk), .Q(ram[3544]) );
  DFFPOSX1 ram_reg_221__7_ ( .D(n7980), .CLK(clk), .Q(ram[3543]) );
  DFFPOSX1 ram_reg_221__6_ ( .D(n7979), .CLK(clk), .Q(ram[3542]) );
  DFFPOSX1 ram_reg_221__5_ ( .D(n7978), .CLK(clk), .Q(ram[3541]) );
  DFFPOSX1 ram_reg_221__4_ ( .D(n7977), .CLK(clk), .Q(ram[3540]) );
  DFFPOSX1 ram_reg_221__3_ ( .D(n7976), .CLK(clk), .Q(ram[3539]) );
  DFFPOSX1 ram_reg_221__2_ ( .D(n7975), .CLK(clk), .Q(ram[3538]) );
  DFFPOSX1 ram_reg_221__1_ ( .D(n7974), .CLK(clk), .Q(ram[3537]) );
  DFFPOSX1 ram_reg_221__0_ ( .D(n7973), .CLK(clk), .Q(ram[3536]) );
  DFFPOSX1 ram_reg_220__15_ ( .D(n7972), .CLK(clk), .Q(ram[3535]) );
  DFFPOSX1 ram_reg_220__14_ ( .D(n7971), .CLK(clk), .Q(ram[3534]) );
  DFFPOSX1 ram_reg_220__13_ ( .D(n7970), .CLK(clk), .Q(ram[3533]) );
  DFFPOSX1 ram_reg_220__12_ ( .D(n7969), .CLK(clk), .Q(ram[3532]) );
  DFFPOSX1 ram_reg_220__11_ ( .D(n7968), .CLK(clk), .Q(ram[3531]) );
  DFFPOSX1 ram_reg_220__10_ ( .D(n7967), .CLK(clk), .Q(ram[3530]) );
  DFFPOSX1 ram_reg_220__9_ ( .D(n7966), .CLK(clk), .Q(ram[3529]) );
  DFFPOSX1 ram_reg_220__8_ ( .D(n7965), .CLK(clk), .Q(ram[3528]) );
  DFFPOSX1 ram_reg_220__7_ ( .D(n7964), .CLK(clk), .Q(ram[3527]) );
  DFFPOSX1 ram_reg_220__6_ ( .D(n7963), .CLK(clk), .Q(ram[3526]) );
  DFFPOSX1 ram_reg_220__5_ ( .D(n7962), .CLK(clk), .Q(ram[3525]) );
  DFFPOSX1 ram_reg_220__4_ ( .D(n7961), .CLK(clk), .Q(ram[3524]) );
  DFFPOSX1 ram_reg_220__3_ ( .D(n7960), .CLK(clk), .Q(ram[3523]) );
  DFFPOSX1 ram_reg_220__2_ ( .D(n7959), .CLK(clk), .Q(ram[3522]) );
  DFFPOSX1 ram_reg_220__1_ ( .D(n7958), .CLK(clk), .Q(ram[3521]) );
  DFFPOSX1 ram_reg_220__0_ ( .D(n7957), .CLK(clk), .Q(ram[3520]) );
  DFFPOSX1 ram_reg_219__15_ ( .D(n7956), .CLK(clk), .Q(ram[3519]) );
  DFFPOSX1 ram_reg_219__14_ ( .D(n7955), .CLK(clk), .Q(ram[3518]) );
  DFFPOSX1 ram_reg_219__13_ ( .D(n7954), .CLK(clk), .Q(ram[3517]) );
  DFFPOSX1 ram_reg_219__12_ ( .D(n7953), .CLK(clk), .Q(ram[3516]) );
  DFFPOSX1 ram_reg_219__11_ ( .D(n7952), .CLK(clk), .Q(ram[3515]) );
  DFFPOSX1 ram_reg_219__10_ ( .D(n7951), .CLK(clk), .Q(ram[3514]) );
  DFFPOSX1 ram_reg_219__9_ ( .D(n7950), .CLK(clk), .Q(ram[3513]) );
  DFFPOSX1 ram_reg_219__8_ ( .D(n7949), .CLK(clk), .Q(ram[3512]) );
  DFFPOSX1 ram_reg_219__7_ ( .D(n7948), .CLK(clk), .Q(ram[3511]) );
  DFFPOSX1 ram_reg_219__6_ ( .D(n7947), .CLK(clk), .Q(ram[3510]) );
  DFFPOSX1 ram_reg_219__5_ ( .D(n7946), .CLK(clk), .Q(ram[3509]) );
  DFFPOSX1 ram_reg_219__4_ ( .D(n7945), .CLK(clk), .Q(ram[3508]) );
  DFFPOSX1 ram_reg_219__3_ ( .D(n7944), .CLK(clk), .Q(ram[3507]) );
  DFFPOSX1 ram_reg_219__2_ ( .D(n7943), .CLK(clk), .Q(ram[3506]) );
  DFFPOSX1 ram_reg_219__1_ ( .D(n7942), .CLK(clk), .Q(ram[3505]) );
  DFFPOSX1 ram_reg_219__0_ ( .D(n7941), .CLK(clk), .Q(ram[3504]) );
  DFFPOSX1 ram_reg_218__15_ ( .D(n7940), .CLK(clk), .Q(ram[3503]) );
  DFFPOSX1 ram_reg_218__14_ ( .D(n7939), .CLK(clk), .Q(ram[3502]) );
  DFFPOSX1 ram_reg_218__13_ ( .D(n7938), .CLK(clk), .Q(ram[3501]) );
  DFFPOSX1 ram_reg_218__12_ ( .D(n7937), .CLK(clk), .Q(ram[3500]) );
  DFFPOSX1 ram_reg_218__11_ ( .D(n7936), .CLK(clk), .Q(ram[3499]) );
  DFFPOSX1 ram_reg_218__10_ ( .D(n7935), .CLK(clk), .Q(ram[3498]) );
  DFFPOSX1 ram_reg_218__9_ ( .D(n7934), .CLK(clk), .Q(ram[3497]) );
  DFFPOSX1 ram_reg_218__8_ ( .D(n7933), .CLK(clk), .Q(ram[3496]) );
  DFFPOSX1 ram_reg_218__7_ ( .D(n7932), .CLK(clk), .Q(ram[3495]) );
  DFFPOSX1 ram_reg_218__6_ ( .D(n7931), .CLK(clk), .Q(ram[3494]) );
  DFFPOSX1 ram_reg_218__5_ ( .D(n7930), .CLK(clk), .Q(ram[3493]) );
  DFFPOSX1 ram_reg_218__4_ ( .D(n7929), .CLK(clk), .Q(ram[3492]) );
  DFFPOSX1 ram_reg_218__3_ ( .D(n7928), .CLK(clk), .Q(ram[3491]) );
  DFFPOSX1 ram_reg_218__2_ ( .D(n7927), .CLK(clk), .Q(ram[3490]) );
  DFFPOSX1 ram_reg_218__1_ ( .D(n7926), .CLK(clk), .Q(ram[3489]) );
  DFFPOSX1 ram_reg_218__0_ ( .D(n7925), .CLK(clk), .Q(ram[3488]) );
  DFFPOSX1 ram_reg_217__15_ ( .D(n7924), .CLK(clk), .Q(ram[3487]) );
  DFFPOSX1 ram_reg_217__14_ ( .D(n7923), .CLK(clk), .Q(ram[3486]) );
  DFFPOSX1 ram_reg_217__13_ ( .D(n7922), .CLK(clk), .Q(ram[3485]) );
  DFFPOSX1 ram_reg_217__12_ ( .D(n7921), .CLK(clk), .Q(ram[3484]) );
  DFFPOSX1 ram_reg_217__11_ ( .D(n7920), .CLK(clk), .Q(ram[3483]) );
  DFFPOSX1 ram_reg_217__10_ ( .D(n7919), .CLK(clk), .Q(ram[3482]) );
  DFFPOSX1 ram_reg_217__9_ ( .D(n7918), .CLK(clk), .Q(ram[3481]) );
  DFFPOSX1 ram_reg_217__8_ ( .D(n7917), .CLK(clk), .Q(ram[3480]) );
  DFFPOSX1 ram_reg_217__7_ ( .D(n7916), .CLK(clk), .Q(ram[3479]) );
  DFFPOSX1 ram_reg_217__6_ ( .D(n7915), .CLK(clk), .Q(ram[3478]) );
  DFFPOSX1 ram_reg_217__5_ ( .D(n7914), .CLK(clk), .Q(ram[3477]) );
  DFFPOSX1 ram_reg_217__4_ ( .D(n7913), .CLK(clk), .Q(ram[3476]) );
  DFFPOSX1 ram_reg_217__3_ ( .D(n7912), .CLK(clk), .Q(ram[3475]) );
  DFFPOSX1 ram_reg_217__2_ ( .D(n7911), .CLK(clk), .Q(ram[3474]) );
  DFFPOSX1 ram_reg_217__1_ ( .D(n7910), .CLK(clk), .Q(ram[3473]) );
  DFFPOSX1 ram_reg_217__0_ ( .D(n7909), .CLK(clk), .Q(ram[3472]) );
  DFFPOSX1 ram_reg_216__15_ ( .D(n7908), .CLK(clk), .Q(ram[3471]) );
  DFFPOSX1 ram_reg_216__14_ ( .D(n7907), .CLK(clk), .Q(ram[3470]) );
  DFFPOSX1 ram_reg_216__13_ ( .D(n7906), .CLK(clk), .Q(ram[3469]) );
  DFFPOSX1 ram_reg_216__12_ ( .D(n7905), .CLK(clk), .Q(ram[3468]) );
  DFFPOSX1 ram_reg_216__11_ ( .D(n7904), .CLK(clk), .Q(ram[3467]) );
  DFFPOSX1 ram_reg_216__10_ ( .D(n7903), .CLK(clk), .Q(ram[3466]) );
  DFFPOSX1 ram_reg_216__9_ ( .D(n7902), .CLK(clk), .Q(ram[3465]) );
  DFFPOSX1 ram_reg_216__8_ ( .D(n7901), .CLK(clk), .Q(ram[3464]) );
  DFFPOSX1 ram_reg_216__7_ ( .D(n7900), .CLK(clk), .Q(ram[3463]) );
  DFFPOSX1 ram_reg_216__6_ ( .D(n7899), .CLK(clk), .Q(ram[3462]) );
  DFFPOSX1 ram_reg_216__5_ ( .D(n7898), .CLK(clk), .Q(ram[3461]) );
  DFFPOSX1 ram_reg_216__4_ ( .D(n7897), .CLK(clk), .Q(ram[3460]) );
  DFFPOSX1 ram_reg_216__3_ ( .D(n7896), .CLK(clk), .Q(ram[3459]) );
  DFFPOSX1 ram_reg_216__2_ ( .D(n7895), .CLK(clk), .Q(ram[3458]) );
  DFFPOSX1 ram_reg_216__1_ ( .D(n7894), .CLK(clk), .Q(ram[3457]) );
  DFFPOSX1 ram_reg_216__0_ ( .D(n7893), .CLK(clk), .Q(ram[3456]) );
  DFFPOSX1 ram_reg_215__15_ ( .D(n7892), .CLK(clk), .Q(ram[3455]) );
  DFFPOSX1 ram_reg_215__14_ ( .D(n7891), .CLK(clk), .Q(ram[3454]) );
  DFFPOSX1 ram_reg_215__13_ ( .D(n7890), .CLK(clk), .Q(ram[3453]) );
  DFFPOSX1 ram_reg_215__12_ ( .D(n7889), .CLK(clk), .Q(ram[3452]) );
  DFFPOSX1 ram_reg_215__11_ ( .D(n7888), .CLK(clk), .Q(ram[3451]) );
  DFFPOSX1 ram_reg_215__10_ ( .D(n7887), .CLK(clk), .Q(ram[3450]) );
  DFFPOSX1 ram_reg_215__9_ ( .D(n7886), .CLK(clk), .Q(ram[3449]) );
  DFFPOSX1 ram_reg_215__8_ ( .D(n7885), .CLK(clk), .Q(ram[3448]) );
  DFFPOSX1 ram_reg_215__7_ ( .D(n7884), .CLK(clk), .Q(ram[3447]) );
  DFFPOSX1 ram_reg_215__6_ ( .D(n7883), .CLK(clk), .Q(ram[3446]) );
  DFFPOSX1 ram_reg_215__5_ ( .D(n7882), .CLK(clk), .Q(ram[3445]) );
  DFFPOSX1 ram_reg_215__4_ ( .D(n7881), .CLK(clk), .Q(ram[3444]) );
  DFFPOSX1 ram_reg_215__3_ ( .D(n7880), .CLK(clk), .Q(ram[3443]) );
  DFFPOSX1 ram_reg_215__2_ ( .D(n7879), .CLK(clk), .Q(ram[3442]) );
  DFFPOSX1 ram_reg_215__1_ ( .D(n7878), .CLK(clk), .Q(ram[3441]) );
  DFFPOSX1 ram_reg_215__0_ ( .D(n7877), .CLK(clk), .Q(ram[3440]) );
  DFFPOSX1 ram_reg_214__15_ ( .D(n7876), .CLK(clk), .Q(ram[3439]) );
  DFFPOSX1 ram_reg_214__14_ ( .D(n7875), .CLK(clk), .Q(ram[3438]) );
  DFFPOSX1 ram_reg_214__13_ ( .D(n7874), .CLK(clk), .Q(ram[3437]) );
  DFFPOSX1 ram_reg_214__12_ ( .D(n7873), .CLK(clk), .Q(ram[3436]) );
  DFFPOSX1 ram_reg_214__11_ ( .D(n7872), .CLK(clk), .Q(ram[3435]) );
  DFFPOSX1 ram_reg_214__10_ ( .D(n7871), .CLK(clk), .Q(ram[3434]) );
  DFFPOSX1 ram_reg_214__9_ ( .D(n7870), .CLK(clk), .Q(ram[3433]) );
  DFFPOSX1 ram_reg_214__8_ ( .D(n7869), .CLK(clk), .Q(ram[3432]) );
  DFFPOSX1 ram_reg_214__7_ ( .D(n7868), .CLK(clk), .Q(ram[3431]) );
  DFFPOSX1 ram_reg_214__6_ ( .D(n7867), .CLK(clk), .Q(ram[3430]) );
  DFFPOSX1 ram_reg_214__5_ ( .D(n7866), .CLK(clk), .Q(ram[3429]) );
  DFFPOSX1 ram_reg_214__4_ ( .D(n7865), .CLK(clk), .Q(ram[3428]) );
  DFFPOSX1 ram_reg_214__3_ ( .D(n7864), .CLK(clk), .Q(ram[3427]) );
  DFFPOSX1 ram_reg_214__2_ ( .D(n7863), .CLK(clk), .Q(ram[3426]) );
  DFFPOSX1 ram_reg_214__1_ ( .D(n7862), .CLK(clk), .Q(ram[3425]) );
  DFFPOSX1 ram_reg_214__0_ ( .D(n7861), .CLK(clk), .Q(ram[3424]) );
  DFFPOSX1 ram_reg_213__15_ ( .D(n7860), .CLK(clk), .Q(ram[3423]) );
  DFFPOSX1 ram_reg_213__14_ ( .D(n7859), .CLK(clk), .Q(ram[3422]) );
  DFFPOSX1 ram_reg_213__13_ ( .D(n7858), .CLK(clk), .Q(ram[3421]) );
  DFFPOSX1 ram_reg_213__12_ ( .D(n7857), .CLK(clk), .Q(ram[3420]) );
  DFFPOSX1 ram_reg_213__11_ ( .D(n7856), .CLK(clk), .Q(ram[3419]) );
  DFFPOSX1 ram_reg_213__10_ ( .D(n7855), .CLK(clk), .Q(ram[3418]) );
  DFFPOSX1 ram_reg_213__9_ ( .D(n7854), .CLK(clk), .Q(ram[3417]) );
  DFFPOSX1 ram_reg_213__8_ ( .D(n7853), .CLK(clk), .Q(ram[3416]) );
  DFFPOSX1 ram_reg_213__7_ ( .D(n7852), .CLK(clk), .Q(ram[3415]) );
  DFFPOSX1 ram_reg_213__6_ ( .D(n7851), .CLK(clk), .Q(ram[3414]) );
  DFFPOSX1 ram_reg_213__5_ ( .D(n7850), .CLK(clk), .Q(ram[3413]) );
  DFFPOSX1 ram_reg_213__4_ ( .D(n7849), .CLK(clk), .Q(ram[3412]) );
  DFFPOSX1 ram_reg_213__3_ ( .D(n7848), .CLK(clk), .Q(ram[3411]) );
  DFFPOSX1 ram_reg_213__2_ ( .D(n7847), .CLK(clk), .Q(ram[3410]) );
  DFFPOSX1 ram_reg_213__1_ ( .D(n7846), .CLK(clk), .Q(ram[3409]) );
  DFFPOSX1 ram_reg_213__0_ ( .D(n7845), .CLK(clk), .Q(ram[3408]) );
  DFFPOSX1 ram_reg_212__15_ ( .D(n7844), .CLK(clk), .Q(ram[3407]) );
  DFFPOSX1 ram_reg_212__14_ ( .D(n7843), .CLK(clk), .Q(ram[3406]) );
  DFFPOSX1 ram_reg_212__13_ ( .D(n7842), .CLK(clk), .Q(ram[3405]) );
  DFFPOSX1 ram_reg_212__12_ ( .D(n7841), .CLK(clk), .Q(ram[3404]) );
  DFFPOSX1 ram_reg_212__11_ ( .D(n7840), .CLK(clk), .Q(ram[3403]) );
  DFFPOSX1 ram_reg_212__10_ ( .D(n7839), .CLK(clk), .Q(ram[3402]) );
  DFFPOSX1 ram_reg_212__9_ ( .D(n7838), .CLK(clk), .Q(ram[3401]) );
  DFFPOSX1 ram_reg_212__8_ ( .D(n7837), .CLK(clk), .Q(ram[3400]) );
  DFFPOSX1 ram_reg_212__7_ ( .D(n7836), .CLK(clk), .Q(ram[3399]) );
  DFFPOSX1 ram_reg_212__6_ ( .D(n7835), .CLK(clk), .Q(ram[3398]) );
  DFFPOSX1 ram_reg_212__5_ ( .D(n7834), .CLK(clk), .Q(ram[3397]) );
  DFFPOSX1 ram_reg_212__4_ ( .D(n7833), .CLK(clk), .Q(ram[3396]) );
  DFFPOSX1 ram_reg_212__3_ ( .D(n7832), .CLK(clk), .Q(ram[3395]) );
  DFFPOSX1 ram_reg_212__2_ ( .D(n7831), .CLK(clk), .Q(ram[3394]) );
  DFFPOSX1 ram_reg_212__1_ ( .D(n7830), .CLK(clk), .Q(ram[3393]) );
  DFFPOSX1 ram_reg_212__0_ ( .D(n7829), .CLK(clk), .Q(ram[3392]) );
  DFFPOSX1 ram_reg_211__15_ ( .D(n7828), .CLK(clk), .Q(ram[3391]) );
  DFFPOSX1 ram_reg_211__14_ ( .D(n7827), .CLK(clk), .Q(ram[3390]) );
  DFFPOSX1 ram_reg_211__13_ ( .D(n7826), .CLK(clk), .Q(ram[3389]) );
  DFFPOSX1 ram_reg_211__12_ ( .D(n7825), .CLK(clk), .Q(ram[3388]) );
  DFFPOSX1 ram_reg_211__11_ ( .D(n7824), .CLK(clk), .Q(ram[3387]) );
  DFFPOSX1 ram_reg_211__10_ ( .D(n7823), .CLK(clk), .Q(ram[3386]) );
  DFFPOSX1 ram_reg_211__9_ ( .D(n7822), .CLK(clk), .Q(ram[3385]) );
  DFFPOSX1 ram_reg_211__8_ ( .D(n7821), .CLK(clk), .Q(ram[3384]) );
  DFFPOSX1 ram_reg_211__7_ ( .D(n7820), .CLK(clk), .Q(ram[3383]) );
  DFFPOSX1 ram_reg_211__6_ ( .D(n7819), .CLK(clk), .Q(ram[3382]) );
  DFFPOSX1 ram_reg_211__5_ ( .D(n7818), .CLK(clk), .Q(ram[3381]) );
  DFFPOSX1 ram_reg_211__4_ ( .D(n7817), .CLK(clk), .Q(ram[3380]) );
  DFFPOSX1 ram_reg_211__3_ ( .D(n7816), .CLK(clk), .Q(ram[3379]) );
  DFFPOSX1 ram_reg_211__2_ ( .D(n7815), .CLK(clk), .Q(ram[3378]) );
  DFFPOSX1 ram_reg_211__1_ ( .D(n7814), .CLK(clk), .Q(ram[3377]) );
  DFFPOSX1 ram_reg_211__0_ ( .D(n7813), .CLK(clk), .Q(ram[3376]) );
  DFFPOSX1 ram_reg_210__15_ ( .D(n7812), .CLK(clk), .Q(ram[3375]) );
  DFFPOSX1 ram_reg_210__14_ ( .D(n7811), .CLK(clk), .Q(ram[3374]) );
  DFFPOSX1 ram_reg_210__13_ ( .D(n7810), .CLK(clk), .Q(ram[3373]) );
  DFFPOSX1 ram_reg_210__12_ ( .D(n7809), .CLK(clk), .Q(ram[3372]) );
  DFFPOSX1 ram_reg_210__11_ ( .D(n7808), .CLK(clk), .Q(ram[3371]) );
  DFFPOSX1 ram_reg_210__10_ ( .D(n7807), .CLK(clk), .Q(ram[3370]) );
  DFFPOSX1 ram_reg_210__9_ ( .D(n7806), .CLK(clk), .Q(ram[3369]) );
  DFFPOSX1 ram_reg_210__8_ ( .D(n7805), .CLK(clk), .Q(ram[3368]) );
  DFFPOSX1 ram_reg_210__7_ ( .D(n7804), .CLK(clk), .Q(ram[3367]) );
  DFFPOSX1 ram_reg_210__6_ ( .D(n7803), .CLK(clk), .Q(ram[3366]) );
  DFFPOSX1 ram_reg_210__5_ ( .D(n7802), .CLK(clk), .Q(ram[3365]) );
  DFFPOSX1 ram_reg_210__4_ ( .D(n7801), .CLK(clk), .Q(ram[3364]) );
  DFFPOSX1 ram_reg_210__3_ ( .D(n7800), .CLK(clk), .Q(ram[3363]) );
  DFFPOSX1 ram_reg_210__2_ ( .D(n7799), .CLK(clk), .Q(ram[3362]) );
  DFFPOSX1 ram_reg_210__1_ ( .D(n7798), .CLK(clk), .Q(ram[3361]) );
  DFFPOSX1 ram_reg_210__0_ ( .D(n7797), .CLK(clk), .Q(ram[3360]) );
  DFFPOSX1 ram_reg_209__15_ ( .D(n7796), .CLK(clk), .Q(ram[3359]) );
  DFFPOSX1 ram_reg_209__14_ ( .D(n7795), .CLK(clk), .Q(ram[3358]) );
  DFFPOSX1 ram_reg_209__13_ ( .D(n7794), .CLK(clk), .Q(ram[3357]) );
  DFFPOSX1 ram_reg_209__12_ ( .D(n7793), .CLK(clk), .Q(ram[3356]) );
  DFFPOSX1 ram_reg_209__11_ ( .D(n7792), .CLK(clk), .Q(ram[3355]) );
  DFFPOSX1 ram_reg_209__10_ ( .D(n7791), .CLK(clk), .Q(ram[3354]) );
  DFFPOSX1 ram_reg_209__9_ ( .D(n7790), .CLK(clk), .Q(ram[3353]) );
  DFFPOSX1 ram_reg_209__8_ ( .D(n7789), .CLK(clk), .Q(ram[3352]) );
  DFFPOSX1 ram_reg_209__7_ ( .D(n7788), .CLK(clk), .Q(ram[3351]) );
  DFFPOSX1 ram_reg_209__6_ ( .D(n7787), .CLK(clk), .Q(ram[3350]) );
  DFFPOSX1 ram_reg_209__5_ ( .D(n7786), .CLK(clk), .Q(ram[3349]) );
  DFFPOSX1 ram_reg_209__4_ ( .D(n7785), .CLK(clk), .Q(ram[3348]) );
  DFFPOSX1 ram_reg_209__3_ ( .D(n7784), .CLK(clk), .Q(ram[3347]) );
  DFFPOSX1 ram_reg_209__2_ ( .D(n7783), .CLK(clk), .Q(ram[3346]) );
  DFFPOSX1 ram_reg_209__1_ ( .D(n7782), .CLK(clk), .Q(ram[3345]) );
  DFFPOSX1 ram_reg_209__0_ ( .D(n7781), .CLK(clk), .Q(ram[3344]) );
  DFFPOSX1 ram_reg_208__15_ ( .D(n7780), .CLK(clk), .Q(ram[3343]) );
  DFFPOSX1 ram_reg_208__14_ ( .D(n7779), .CLK(clk), .Q(ram[3342]) );
  DFFPOSX1 ram_reg_208__13_ ( .D(n7778), .CLK(clk), .Q(ram[3341]) );
  DFFPOSX1 ram_reg_208__12_ ( .D(n7777), .CLK(clk), .Q(ram[3340]) );
  DFFPOSX1 ram_reg_208__11_ ( .D(n7776), .CLK(clk), .Q(ram[3339]) );
  DFFPOSX1 ram_reg_208__10_ ( .D(n7775), .CLK(clk), .Q(ram[3338]) );
  DFFPOSX1 ram_reg_208__9_ ( .D(n7774), .CLK(clk), .Q(ram[3337]) );
  DFFPOSX1 ram_reg_208__8_ ( .D(n7773), .CLK(clk), .Q(ram[3336]) );
  DFFPOSX1 ram_reg_208__7_ ( .D(n7772), .CLK(clk), .Q(ram[3335]) );
  DFFPOSX1 ram_reg_208__6_ ( .D(n7771), .CLK(clk), .Q(ram[3334]) );
  DFFPOSX1 ram_reg_208__5_ ( .D(n7770), .CLK(clk), .Q(ram[3333]) );
  DFFPOSX1 ram_reg_208__4_ ( .D(n7769), .CLK(clk), .Q(ram[3332]) );
  DFFPOSX1 ram_reg_208__3_ ( .D(n7768), .CLK(clk), .Q(ram[3331]) );
  DFFPOSX1 ram_reg_208__2_ ( .D(n7767), .CLK(clk), .Q(ram[3330]) );
  DFFPOSX1 ram_reg_208__1_ ( .D(n7766), .CLK(clk), .Q(ram[3329]) );
  DFFPOSX1 ram_reg_208__0_ ( .D(n7765), .CLK(clk), .Q(ram[3328]) );
  DFFPOSX1 ram_reg_207__15_ ( .D(n7764), .CLK(clk), .Q(ram[3327]) );
  DFFPOSX1 ram_reg_207__14_ ( .D(n7763), .CLK(clk), .Q(ram[3326]) );
  DFFPOSX1 ram_reg_207__13_ ( .D(n7762), .CLK(clk), .Q(ram[3325]) );
  DFFPOSX1 ram_reg_207__12_ ( .D(n7761), .CLK(clk), .Q(ram[3324]) );
  DFFPOSX1 ram_reg_207__11_ ( .D(n7760), .CLK(clk), .Q(ram[3323]) );
  DFFPOSX1 ram_reg_207__10_ ( .D(n7759), .CLK(clk), .Q(ram[3322]) );
  DFFPOSX1 ram_reg_207__9_ ( .D(n7758), .CLK(clk), .Q(ram[3321]) );
  DFFPOSX1 ram_reg_207__8_ ( .D(n7757), .CLK(clk), .Q(ram[3320]) );
  DFFPOSX1 ram_reg_207__7_ ( .D(n7756), .CLK(clk), .Q(ram[3319]) );
  DFFPOSX1 ram_reg_207__6_ ( .D(n7755), .CLK(clk), .Q(ram[3318]) );
  DFFPOSX1 ram_reg_207__5_ ( .D(n7754), .CLK(clk), .Q(ram[3317]) );
  DFFPOSX1 ram_reg_207__4_ ( .D(n7753), .CLK(clk), .Q(ram[3316]) );
  DFFPOSX1 ram_reg_207__3_ ( .D(n7752), .CLK(clk), .Q(ram[3315]) );
  DFFPOSX1 ram_reg_207__2_ ( .D(n7751), .CLK(clk), .Q(ram[3314]) );
  DFFPOSX1 ram_reg_207__1_ ( .D(n7750), .CLK(clk), .Q(ram[3313]) );
  DFFPOSX1 ram_reg_207__0_ ( .D(n7749), .CLK(clk), .Q(ram[3312]) );
  DFFPOSX1 ram_reg_206__15_ ( .D(n7748), .CLK(clk), .Q(ram[3311]) );
  DFFPOSX1 ram_reg_206__14_ ( .D(n7747), .CLK(clk), .Q(ram[3310]) );
  DFFPOSX1 ram_reg_206__13_ ( .D(n7746), .CLK(clk), .Q(ram[3309]) );
  DFFPOSX1 ram_reg_206__12_ ( .D(n7745), .CLK(clk), .Q(ram[3308]) );
  DFFPOSX1 ram_reg_206__11_ ( .D(n7744), .CLK(clk), .Q(ram[3307]) );
  DFFPOSX1 ram_reg_206__10_ ( .D(n7743), .CLK(clk), .Q(ram[3306]) );
  DFFPOSX1 ram_reg_206__9_ ( .D(n7742), .CLK(clk), .Q(ram[3305]) );
  DFFPOSX1 ram_reg_206__8_ ( .D(n7741), .CLK(clk), .Q(ram[3304]) );
  DFFPOSX1 ram_reg_206__7_ ( .D(n7740), .CLK(clk), .Q(ram[3303]) );
  DFFPOSX1 ram_reg_206__6_ ( .D(n7739), .CLK(clk), .Q(ram[3302]) );
  DFFPOSX1 ram_reg_206__5_ ( .D(n7738), .CLK(clk), .Q(ram[3301]) );
  DFFPOSX1 ram_reg_206__4_ ( .D(n7737), .CLK(clk), .Q(ram[3300]) );
  DFFPOSX1 ram_reg_206__3_ ( .D(n7736), .CLK(clk), .Q(ram[3299]) );
  DFFPOSX1 ram_reg_206__2_ ( .D(n7735), .CLK(clk), .Q(ram[3298]) );
  DFFPOSX1 ram_reg_206__1_ ( .D(n7734), .CLK(clk), .Q(ram[3297]) );
  DFFPOSX1 ram_reg_206__0_ ( .D(n7733), .CLK(clk), .Q(ram[3296]) );
  DFFPOSX1 ram_reg_205__15_ ( .D(n7732), .CLK(clk), .Q(ram[3295]) );
  DFFPOSX1 ram_reg_205__14_ ( .D(n7731), .CLK(clk), .Q(ram[3294]) );
  DFFPOSX1 ram_reg_205__13_ ( .D(n7730), .CLK(clk), .Q(ram[3293]) );
  DFFPOSX1 ram_reg_205__12_ ( .D(n7729), .CLK(clk), .Q(ram[3292]) );
  DFFPOSX1 ram_reg_205__11_ ( .D(n7728), .CLK(clk), .Q(ram[3291]) );
  DFFPOSX1 ram_reg_205__10_ ( .D(n7727), .CLK(clk), .Q(ram[3290]) );
  DFFPOSX1 ram_reg_205__9_ ( .D(n7726), .CLK(clk), .Q(ram[3289]) );
  DFFPOSX1 ram_reg_205__8_ ( .D(n7725), .CLK(clk), .Q(ram[3288]) );
  DFFPOSX1 ram_reg_205__7_ ( .D(n7724), .CLK(clk), .Q(ram[3287]) );
  DFFPOSX1 ram_reg_205__6_ ( .D(n7723), .CLK(clk), .Q(ram[3286]) );
  DFFPOSX1 ram_reg_205__5_ ( .D(n7722), .CLK(clk), .Q(ram[3285]) );
  DFFPOSX1 ram_reg_205__4_ ( .D(n7721), .CLK(clk), .Q(ram[3284]) );
  DFFPOSX1 ram_reg_205__3_ ( .D(n7720), .CLK(clk), .Q(ram[3283]) );
  DFFPOSX1 ram_reg_205__2_ ( .D(n7719), .CLK(clk), .Q(ram[3282]) );
  DFFPOSX1 ram_reg_205__1_ ( .D(n7718), .CLK(clk), .Q(ram[3281]) );
  DFFPOSX1 ram_reg_205__0_ ( .D(n7717), .CLK(clk), .Q(ram[3280]) );
  DFFPOSX1 ram_reg_204__15_ ( .D(n7716), .CLK(clk), .Q(ram[3279]) );
  DFFPOSX1 ram_reg_204__14_ ( .D(n7715), .CLK(clk), .Q(ram[3278]) );
  DFFPOSX1 ram_reg_204__13_ ( .D(n7714), .CLK(clk), .Q(ram[3277]) );
  DFFPOSX1 ram_reg_204__12_ ( .D(n7713), .CLK(clk), .Q(ram[3276]) );
  DFFPOSX1 ram_reg_204__11_ ( .D(n7712), .CLK(clk), .Q(ram[3275]) );
  DFFPOSX1 ram_reg_204__10_ ( .D(n7711), .CLK(clk), .Q(ram[3274]) );
  DFFPOSX1 ram_reg_204__9_ ( .D(n7710), .CLK(clk), .Q(ram[3273]) );
  DFFPOSX1 ram_reg_204__8_ ( .D(n7709), .CLK(clk), .Q(ram[3272]) );
  DFFPOSX1 ram_reg_204__7_ ( .D(n7708), .CLK(clk), .Q(ram[3271]) );
  DFFPOSX1 ram_reg_204__6_ ( .D(n7707), .CLK(clk), .Q(ram[3270]) );
  DFFPOSX1 ram_reg_204__5_ ( .D(n7706), .CLK(clk), .Q(ram[3269]) );
  DFFPOSX1 ram_reg_204__4_ ( .D(n7705), .CLK(clk), .Q(ram[3268]) );
  DFFPOSX1 ram_reg_204__3_ ( .D(n7704), .CLK(clk), .Q(ram[3267]) );
  DFFPOSX1 ram_reg_204__2_ ( .D(n7703), .CLK(clk), .Q(ram[3266]) );
  DFFPOSX1 ram_reg_204__1_ ( .D(n7702), .CLK(clk), .Q(ram[3265]) );
  DFFPOSX1 ram_reg_204__0_ ( .D(n7701), .CLK(clk), .Q(ram[3264]) );
  DFFPOSX1 ram_reg_203__15_ ( .D(n7700), .CLK(clk), .Q(ram[3263]) );
  DFFPOSX1 ram_reg_203__14_ ( .D(n7699), .CLK(clk), .Q(ram[3262]) );
  DFFPOSX1 ram_reg_203__13_ ( .D(n7698), .CLK(clk), .Q(ram[3261]) );
  DFFPOSX1 ram_reg_203__12_ ( .D(n7697), .CLK(clk), .Q(ram[3260]) );
  DFFPOSX1 ram_reg_203__11_ ( .D(n7696), .CLK(clk), .Q(ram[3259]) );
  DFFPOSX1 ram_reg_203__10_ ( .D(n7695), .CLK(clk), .Q(ram[3258]) );
  DFFPOSX1 ram_reg_203__9_ ( .D(n7694), .CLK(clk), .Q(ram[3257]) );
  DFFPOSX1 ram_reg_203__8_ ( .D(n7693), .CLK(clk), .Q(ram[3256]) );
  DFFPOSX1 ram_reg_203__7_ ( .D(n7692), .CLK(clk), .Q(ram[3255]) );
  DFFPOSX1 ram_reg_203__6_ ( .D(n7691), .CLK(clk), .Q(ram[3254]) );
  DFFPOSX1 ram_reg_203__5_ ( .D(n7690), .CLK(clk), .Q(ram[3253]) );
  DFFPOSX1 ram_reg_203__4_ ( .D(n7689), .CLK(clk), .Q(ram[3252]) );
  DFFPOSX1 ram_reg_203__3_ ( .D(n7688), .CLK(clk), .Q(ram[3251]) );
  DFFPOSX1 ram_reg_203__2_ ( .D(n7687), .CLK(clk), .Q(ram[3250]) );
  DFFPOSX1 ram_reg_203__1_ ( .D(n7686), .CLK(clk), .Q(ram[3249]) );
  DFFPOSX1 ram_reg_203__0_ ( .D(n7685), .CLK(clk), .Q(ram[3248]) );
  DFFPOSX1 ram_reg_202__15_ ( .D(n7684), .CLK(clk), .Q(ram[3247]) );
  DFFPOSX1 ram_reg_202__14_ ( .D(n7683), .CLK(clk), .Q(ram[3246]) );
  DFFPOSX1 ram_reg_202__13_ ( .D(n7682), .CLK(clk), .Q(ram[3245]) );
  DFFPOSX1 ram_reg_202__12_ ( .D(n7681), .CLK(clk), .Q(ram[3244]) );
  DFFPOSX1 ram_reg_202__11_ ( .D(n7680), .CLK(clk), .Q(ram[3243]) );
  DFFPOSX1 ram_reg_202__10_ ( .D(n7679), .CLK(clk), .Q(ram[3242]) );
  DFFPOSX1 ram_reg_202__9_ ( .D(n7678), .CLK(clk), .Q(ram[3241]) );
  DFFPOSX1 ram_reg_202__8_ ( .D(n7677), .CLK(clk), .Q(ram[3240]) );
  DFFPOSX1 ram_reg_202__7_ ( .D(n7676), .CLK(clk), .Q(ram[3239]) );
  DFFPOSX1 ram_reg_202__6_ ( .D(n7675), .CLK(clk), .Q(ram[3238]) );
  DFFPOSX1 ram_reg_202__5_ ( .D(n7674), .CLK(clk), .Q(ram[3237]) );
  DFFPOSX1 ram_reg_202__4_ ( .D(n7673), .CLK(clk), .Q(ram[3236]) );
  DFFPOSX1 ram_reg_202__3_ ( .D(n7672), .CLK(clk), .Q(ram[3235]) );
  DFFPOSX1 ram_reg_202__2_ ( .D(n7671), .CLK(clk), .Q(ram[3234]) );
  DFFPOSX1 ram_reg_202__1_ ( .D(n7670), .CLK(clk), .Q(ram[3233]) );
  DFFPOSX1 ram_reg_202__0_ ( .D(n7669), .CLK(clk), .Q(ram[3232]) );
  DFFPOSX1 ram_reg_201__15_ ( .D(n7668), .CLK(clk), .Q(ram[3231]) );
  DFFPOSX1 ram_reg_201__14_ ( .D(n7667), .CLK(clk), .Q(ram[3230]) );
  DFFPOSX1 ram_reg_201__13_ ( .D(n7666), .CLK(clk), .Q(ram[3229]) );
  DFFPOSX1 ram_reg_201__12_ ( .D(n7665), .CLK(clk), .Q(ram[3228]) );
  DFFPOSX1 ram_reg_201__11_ ( .D(n7664), .CLK(clk), .Q(ram[3227]) );
  DFFPOSX1 ram_reg_201__10_ ( .D(n7663), .CLK(clk), .Q(ram[3226]) );
  DFFPOSX1 ram_reg_201__9_ ( .D(n7662), .CLK(clk), .Q(ram[3225]) );
  DFFPOSX1 ram_reg_201__8_ ( .D(n7661), .CLK(clk), .Q(ram[3224]) );
  DFFPOSX1 ram_reg_201__7_ ( .D(n7660), .CLK(clk), .Q(ram[3223]) );
  DFFPOSX1 ram_reg_201__6_ ( .D(n7659), .CLK(clk), .Q(ram[3222]) );
  DFFPOSX1 ram_reg_201__5_ ( .D(n7658), .CLK(clk), .Q(ram[3221]) );
  DFFPOSX1 ram_reg_201__4_ ( .D(n7657), .CLK(clk), .Q(ram[3220]) );
  DFFPOSX1 ram_reg_201__3_ ( .D(n7656), .CLK(clk), .Q(ram[3219]) );
  DFFPOSX1 ram_reg_201__2_ ( .D(n7655), .CLK(clk), .Q(ram[3218]) );
  DFFPOSX1 ram_reg_201__1_ ( .D(n7654), .CLK(clk), .Q(ram[3217]) );
  DFFPOSX1 ram_reg_201__0_ ( .D(n7653), .CLK(clk), .Q(ram[3216]) );
  DFFPOSX1 ram_reg_200__15_ ( .D(n7652), .CLK(clk), .Q(ram[3215]) );
  DFFPOSX1 ram_reg_200__14_ ( .D(n7651), .CLK(clk), .Q(ram[3214]) );
  DFFPOSX1 ram_reg_200__13_ ( .D(n7650), .CLK(clk), .Q(ram[3213]) );
  DFFPOSX1 ram_reg_200__12_ ( .D(n7649), .CLK(clk), .Q(ram[3212]) );
  DFFPOSX1 ram_reg_200__11_ ( .D(n7648), .CLK(clk), .Q(ram[3211]) );
  DFFPOSX1 ram_reg_200__10_ ( .D(n7647), .CLK(clk), .Q(ram[3210]) );
  DFFPOSX1 ram_reg_200__9_ ( .D(n7646), .CLK(clk), .Q(ram[3209]) );
  DFFPOSX1 ram_reg_200__8_ ( .D(n7645), .CLK(clk), .Q(ram[3208]) );
  DFFPOSX1 ram_reg_200__7_ ( .D(n7644), .CLK(clk), .Q(ram[3207]) );
  DFFPOSX1 ram_reg_200__6_ ( .D(n7643), .CLK(clk), .Q(ram[3206]) );
  DFFPOSX1 ram_reg_200__5_ ( .D(n7642), .CLK(clk), .Q(ram[3205]) );
  DFFPOSX1 ram_reg_200__4_ ( .D(n7641), .CLK(clk), .Q(ram[3204]) );
  DFFPOSX1 ram_reg_200__3_ ( .D(n7640), .CLK(clk), .Q(ram[3203]) );
  DFFPOSX1 ram_reg_200__2_ ( .D(n7639), .CLK(clk), .Q(ram[3202]) );
  DFFPOSX1 ram_reg_200__1_ ( .D(n7638), .CLK(clk), .Q(ram[3201]) );
  DFFPOSX1 ram_reg_200__0_ ( .D(n7637), .CLK(clk), .Q(ram[3200]) );
  DFFPOSX1 ram_reg_199__15_ ( .D(n7636), .CLK(clk), .Q(ram[3199]) );
  DFFPOSX1 ram_reg_199__14_ ( .D(n7635), .CLK(clk), .Q(ram[3198]) );
  DFFPOSX1 ram_reg_199__13_ ( .D(n7634), .CLK(clk), .Q(ram[3197]) );
  DFFPOSX1 ram_reg_199__12_ ( .D(n7633), .CLK(clk), .Q(ram[3196]) );
  DFFPOSX1 ram_reg_199__11_ ( .D(n7632), .CLK(clk), .Q(ram[3195]) );
  DFFPOSX1 ram_reg_199__10_ ( .D(n7631), .CLK(clk), .Q(ram[3194]) );
  DFFPOSX1 ram_reg_199__9_ ( .D(n7630), .CLK(clk), .Q(ram[3193]) );
  DFFPOSX1 ram_reg_199__8_ ( .D(n7629), .CLK(clk), .Q(ram[3192]) );
  DFFPOSX1 ram_reg_199__7_ ( .D(n7628), .CLK(clk), .Q(ram[3191]) );
  DFFPOSX1 ram_reg_199__6_ ( .D(n7627), .CLK(clk), .Q(ram[3190]) );
  DFFPOSX1 ram_reg_199__5_ ( .D(n7626), .CLK(clk), .Q(ram[3189]) );
  DFFPOSX1 ram_reg_199__4_ ( .D(n7625), .CLK(clk), .Q(ram[3188]) );
  DFFPOSX1 ram_reg_199__3_ ( .D(n7624), .CLK(clk), .Q(ram[3187]) );
  DFFPOSX1 ram_reg_199__2_ ( .D(n7623), .CLK(clk), .Q(ram[3186]) );
  DFFPOSX1 ram_reg_199__1_ ( .D(n7622), .CLK(clk), .Q(ram[3185]) );
  DFFPOSX1 ram_reg_199__0_ ( .D(n7621), .CLK(clk), .Q(ram[3184]) );
  DFFPOSX1 ram_reg_198__15_ ( .D(n7620), .CLK(clk), .Q(ram[3183]) );
  DFFPOSX1 ram_reg_198__14_ ( .D(n7619), .CLK(clk), .Q(ram[3182]) );
  DFFPOSX1 ram_reg_198__13_ ( .D(n7618), .CLK(clk), .Q(ram[3181]) );
  DFFPOSX1 ram_reg_198__12_ ( .D(n7617), .CLK(clk), .Q(ram[3180]) );
  DFFPOSX1 ram_reg_198__11_ ( .D(n7616), .CLK(clk), .Q(ram[3179]) );
  DFFPOSX1 ram_reg_198__10_ ( .D(n7615), .CLK(clk), .Q(ram[3178]) );
  DFFPOSX1 ram_reg_198__9_ ( .D(n7614), .CLK(clk), .Q(ram[3177]) );
  DFFPOSX1 ram_reg_198__8_ ( .D(n7613), .CLK(clk), .Q(ram[3176]) );
  DFFPOSX1 ram_reg_198__7_ ( .D(n7612), .CLK(clk), .Q(ram[3175]) );
  DFFPOSX1 ram_reg_198__6_ ( .D(n7611), .CLK(clk), .Q(ram[3174]) );
  DFFPOSX1 ram_reg_198__5_ ( .D(n7610), .CLK(clk), .Q(ram[3173]) );
  DFFPOSX1 ram_reg_198__4_ ( .D(n7609), .CLK(clk), .Q(ram[3172]) );
  DFFPOSX1 ram_reg_198__3_ ( .D(n7608), .CLK(clk), .Q(ram[3171]) );
  DFFPOSX1 ram_reg_198__2_ ( .D(n7607), .CLK(clk), .Q(ram[3170]) );
  DFFPOSX1 ram_reg_198__1_ ( .D(n7606), .CLK(clk), .Q(ram[3169]) );
  DFFPOSX1 ram_reg_198__0_ ( .D(n7605), .CLK(clk), .Q(ram[3168]) );
  DFFPOSX1 ram_reg_197__15_ ( .D(n7604), .CLK(clk), .Q(ram[3167]) );
  DFFPOSX1 ram_reg_197__14_ ( .D(n7603), .CLK(clk), .Q(ram[3166]) );
  DFFPOSX1 ram_reg_197__13_ ( .D(n7602), .CLK(clk), .Q(ram[3165]) );
  DFFPOSX1 ram_reg_197__12_ ( .D(n7601), .CLK(clk), .Q(ram[3164]) );
  DFFPOSX1 ram_reg_197__11_ ( .D(n7600), .CLK(clk), .Q(ram[3163]) );
  DFFPOSX1 ram_reg_197__10_ ( .D(n7599), .CLK(clk), .Q(ram[3162]) );
  DFFPOSX1 ram_reg_197__9_ ( .D(n7598), .CLK(clk), .Q(ram[3161]) );
  DFFPOSX1 ram_reg_197__8_ ( .D(n7597), .CLK(clk), .Q(ram[3160]) );
  DFFPOSX1 ram_reg_197__7_ ( .D(n7596), .CLK(clk), .Q(ram[3159]) );
  DFFPOSX1 ram_reg_197__6_ ( .D(n7595), .CLK(clk), .Q(ram[3158]) );
  DFFPOSX1 ram_reg_197__5_ ( .D(n7594), .CLK(clk), .Q(ram[3157]) );
  DFFPOSX1 ram_reg_197__4_ ( .D(n7593), .CLK(clk), .Q(ram[3156]) );
  DFFPOSX1 ram_reg_197__3_ ( .D(n7592), .CLK(clk), .Q(ram[3155]) );
  DFFPOSX1 ram_reg_197__2_ ( .D(n7591), .CLK(clk), .Q(ram[3154]) );
  DFFPOSX1 ram_reg_197__1_ ( .D(n7590), .CLK(clk), .Q(ram[3153]) );
  DFFPOSX1 ram_reg_197__0_ ( .D(n7589), .CLK(clk), .Q(ram[3152]) );
  DFFPOSX1 ram_reg_196__15_ ( .D(n7588), .CLK(clk), .Q(ram[3151]) );
  DFFPOSX1 ram_reg_196__14_ ( .D(n7587), .CLK(clk), .Q(ram[3150]) );
  DFFPOSX1 ram_reg_196__13_ ( .D(n7586), .CLK(clk), .Q(ram[3149]) );
  DFFPOSX1 ram_reg_196__12_ ( .D(n7585), .CLK(clk), .Q(ram[3148]) );
  DFFPOSX1 ram_reg_196__11_ ( .D(n7584), .CLK(clk), .Q(ram[3147]) );
  DFFPOSX1 ram_reg_196__10_ ( .D(n7583), .CLK(clk), .Q(ram[3146]) );
  DFFPOSX1 ram_reg_196__9_ ( .D(n7582), .CLK(clk), .Q(ram[3145]) );
  DFFPOSX1 ram_reg_196__8_ ( .D(n7581), .CLK(clk), .Q(ram[3144]) );
  DFFPOSX1 ram_reg_196__7_ ( .D(n7580), .CLK(clk), .Q(ram[3143]) );
  DFFPOSX1 ram_reg_196__6_ ( .D(n7579), .CLK(clk), .Q(ram[3142]) );
  DFFPOSX1 ram_reg_196__5_ ( .D(n7578), .CLK(clk), .Q(ram[3141]) );
  DFFPOSX1 ram_reg_196__4_ ( .D(n7577), .CLK(clk), .Q(ram[3140]) );
  DFFPOSX1 ram_reg_196__3_ ( .D(n7576), .CLK(clk), .Q(ram[3139]) );
  DFFPOSX1 ram_reg_196__2_ ( .D(n7575), .CLK(clk), .Q(ram[3138]) );
  DFFPOSX1 ram_reg_196__1_ ( .D(n7574), .CLK(clk), .Q(ram[3137]) );
  DFFPOSX1 ram_reg_196__0_ ( .D(n7573), .CLK(clk), .Q(ram[3136]) );
  DFFPOSX1 ram_reg_195__15_ ( .D(n7572), .CLK(clk), .Q(ram[3135]) );
  DFFPOSX1 ram_reg_195__14_ ( .D(n7571), .CLK(clk), .Q(ram[3134]) );
  DFFPOSX1 ram_reg_195__13_ ( .D(n7570), .CLK(clk), .Q(ram[3133]) );
  DFFPOSX1 ram_reg_195__12_ ( .D(n7569), .CLK(clk), .Q(ram[3132]) );
  DFFPOSX1 ram_reg_195__11_ ( .D(n7568), .CLK(clk), .Q(ram[3131]) );
  DFFPOSX1 ram_reg_195__10_ ( .D(n7567), .CLK(clk), .Q(ram[3130]) );
  DFFPOSX1 ram_reg_195__9_ ( .D(n7566), .CLK(clk), .Q(ram[3129]) );
  DFFPOSX1 ram_reg_195__8_ ( .D(n7565), .CLK(clk), .Q(ram[3128]) );
  DFFPOSX1 ram_reg_195__7_ ( .D(n7564), .CLK(clk), .Q(ram[3127]) );
  DFFPOSX1 ram_reg_195__6_ ( .D(n7563), .CLK(clk), .Q(ram[3126]) );
  DFFPOSX1 ram_reg_195__5_ ( .D(n7562), .CLK(clk), .Q(ram[3125]) );
  DFFPOSX1 ram_reg_195__4_ ( .D(n7561), .CLK(clk), .Q(ram[3124]) );
  DFFPOSX1 ram_reg_195__3_ ( .D(n7560), .CLK(clk), .Q(ram[3123]) );
  DFFPOSX1 ram_reg_195__2_ ( .D(n7559), .CLK(clk), .Q(ram[3122]) );
  DFFPOSX1 ram_reg_195__1_ ( .D(n7558), .CLK(clk), .Q(ram[3121]) );
  DFFPOSX1 ram_reg_195__0_ ( .D(n7557), .CLK(clk), .Q(ram[3120]) );
  DFFPOSX1 ram_reg_194__15_ ( .D(n7556), .CLK(clk), .Q(ram[3119]) );
  DFFPOSX1 ram_reg_194__14_ ( .D(n7555), .CLK(clk), .Q(ram[3118]) );
  DFFPOSX1 ram_reg_194__13_ ( .D(n7554), .CLK(clk), .Q(ram[3117]) );
  DFFPOSX1 ram_reg_194__12_ ( .D(n7553), .CLK(clk), .Q(ram[3116]) );
  DFFPOSX1 ram_reg_194__11_ ( .D(n7552), .CLK(clk), .Q(ram[3115]) );
  DFFPOSX1 ram_reg_194__10_ ( .D(n7551), .CLK(clk), .Q(ram[3114]) );
  DFFPOSX1 ram_reg_194__9_ ( .D(n7550), .CLK(clk), .Q(ram[3113]) );
  DFFPOSX1 ram_reg_194__8_ ( .D(n7549), .CLK(clk), .Q(ram[3112]) );
  DFFPOSX1 ram_reg_194__7_ ( .D(n7548), .CLK(clk), .Q(ram[3111]) );
  DFFPOSX1 ram_reg_194__6_ ( .D(n7547), .CLK(clk), .Q(ram[3110]) );
  DFFPOSX1 ram_reg_194__5_ ( .D(n7546), .CLK(clk), .Q(ram[3109]) );
  DFFPOSX1 ram_reg_194__4_ ( .D(n7545), .CLK(clk), .Q(ram[3108]) );
  DFFPOSX1 ram_reg_194__3_ ( .D(n7544), .CLK(clk), .Q(ram[3107]) );
  DFFPOSX1 ram_reg_194__2_ ( .D(n7543), .CLK(clk), .Q(ram[3106]) );
  DFFPOSX1 ram_reg_194__1_ ( .D(n7542), .CLK(clk), .Q(ram[3105]) );
  DFFPOSX1 ram_reg_194__0_ ( .D(n7541), .CLK(clk), .Q(ram[3104]) );
  DFFPOSX1 ram_reg_193__15_ ( .D(n7540), .CLK(clk), .Q(ram[3103]) );
  DFFPOSX1 ram_reg_193__14_ ( .D(n7539), .CLK(clk), .Q(ram[3102]) );
  DFFPOSX1 ram_reg_193__13_ ( .D(n7538), .CLK(clk), .Q(ram[3101]) );
  DFFPOSX1 ram_reg_193__12_ ( .D(n7537), .CLK(clk), .Q(ram[3100]) );
  DFFPOSX1 ram_reg_193__11_ ( .D(n7536), .CLK(clk), .Q(ram[3099]) );
  DFFPOSX1 ram_reg_193__10_ ( .D(n7535), .CLK(clk), .Q(ram[3098]) );
  DFFPOSX1 ram_reg_193__9_ ( .D(n7534), .CLK(clk), .Q(ram[3097]) );
  DFFPOSX1 ram_reg_193__8_ ( .D(n7533), .CLK(clk), .Q(ram[3096]) );
  DFFPOSX1 ram_reg_193__7_ ( .D(n7532), .CLK(clk), .Q(ram[3095]) );
  DFFPOSX1 ram_reg_193__6_ ( .D(n7531), .CLK(clk), .Q(ram[3094]) );
  DFFPOSX1 ram_reg_193__5_ ( .D(n7530), .CLK(clk), .Q(ram[3093]) );
  DFFPOSX1 ram_reg_193__4_ ( .D(n7529), .CLK(clk), .Q(ram[3092]) );
  DFFPOSX1 ram_reg_193__3_ ( .D(n7528), .CLK(clk), .Q(ram[3091]) );
  DFFPOSX1 ram_reg_193__2_ ( .D(n7527), .CLK(clk), .Q(ram[3090]) );
  DFFPOSX1 ram_reg_193__1_ ( .D(n7526), .CLK(clk), .Q(ram[3089]) );
  DFFPOSX1 ram_reg_193__0_ ( .D(n7525), .CLK(clk), .Q(ram[3088]) );
  DFFPOSX1 ram_reg_192__15_ ( .D(n7524), .CLK(clk), .Q(ram[3087]) );
  DFFPOSX1 ram_reg_192__14_ ( .D(n7523), .CLK(clk), .Q(ram[3086]) );
  DFFPOSX1 ram_reg_192__13_ ( .D(n7522), .CLK(clk), .Q(ram[3085]) );
  DFFPOSX1 ram_reg_192__12_ ( .D(n7521), .CLK(clk), .Q(ram[3084]) );
  DFFPOSX1 ram_reg_192__11_ ( .D(n7520), .CLK(clk), .Q(ram[3083]) );
  DFFPOSX1 ram_reg_192__10_ ( .D(n7519), .CLK(clk), .Q(ram[3082]) );
  DFFPOSX1 ram_reg_192__9_ ( .D(n7518), .CLK(clk), .Q(ram[3081]) );
  DFFPOSX1 ram_reg_192__8_ ( .D(n7517), .CLK(clk), .Q(ram[3080]) );
  DFFPOSX1 ram_reg_192__7_ ( .D(n7516), .CLK(clk), .Q(ram[3079]) );
  DFFPOSX1 ram_reg_192__6_ ( .D(n7515), .CLK(clk), .Q(ram[3078]) );
  DFFPOSX1 ram_reg_192__5_ ( .D(n7514), .CLK(clk), .Q(ram[3077]) );
  DFFPOSX1 ram_reg_192__4_ ( .D(n7513), .CLK(clk), .Q(ram[3076]) );
  DFFPOSX1 ram_reg_192__3_ ( .D(n7512), .CLK(clk), .Q(ram[3075]) );
  DFFPOSX1 ram_reg_192__2_ ( .D(n7511), .CLK(clk), .Q(ram[3074]) );
  DFFPOSX1 ram_reg_192__1_ ( .D(n7510), .CLK(clk), .Q(ram[3073]) );
  DFFPOSX1 ram_reg_192__0_ ( .D(n7509), .CLK(clk), .Q(ram[3072]) );
  DFFPOSX1 ram_reg_191__15_ ( .D(n7508), .CLK(clk), .Q(ram[3071]) );
  DFFPOSX1 ram_reg_191__14_ ( .D(n7507), .CLK(clk), .Q(ram[3070]) );
  DFFPOSX1 ram_reg_191__13_ ( .D(n7506), .CLK(clk), .Q(ram[3069]) );
  DFFPOSX1 ram_reg_191__12_ ( .D(n7505), .CLK(clk), .Q(ram[3068]) );
  DFFPOSX1 ram_reg_191__11_ ( .D(n7504), .CLK(clk), .Q(ram[3067]) );
  DFFPOSX1 ram_reg_191__10_ ( .D(n7503), .CLK(clk), .Q(ram[3066]) );
  DFFPOSX1 ram_reg_191__9_ ( .D(n7502), .CLK(clk), .Q(ram[3065]) );
  DFFPOSX1 ram_reg_191__8_ ( .D(n7501), .CLK(clk), .Q(ram[3064]) );
  DFFPOSX1 ram_reg_191__7_ ( .D(n7500), .CLK(clk), .Q(ram[3063]) );
  DFFPOSX1 ram_reg_191__6_ ( .D(n7499), .CLK(clk), .Q(ram[3062]) );
  DFFPOSX1 ram_reg_191__5_ ( .D(n7498), .CLK(clk), .Q(ram[3061]) );
  DFFPOSX1 ram_reg_191__4_ ( .D(n7497), .CLK(clk), .Q(ram[3060]) );
  DFFPOSX1 ram_reg_191__3_ ( .D(n7496), .CLK(clk), .Q(ram[3059]) );
  DFFPOSX1 ram_reg_191__2_ ( .D(n7495), .CLK(clk), .Q(ram[3058]) );
  DFFPOSX1 ram_reg_191__1_ ( .D(n7494), .CLK(clk), .Q(ram[3057]) );
  DFFPOSX1 ram_reg_191__0_ ( .D(n7493), .CLK(clk), .Q(ram[3056]) );
  DFFPOSX1 ram_reg_190__15_ ( .D(n7492), .CLK(clk), .Q(ram[3055]) );
  DFFPOSX1 ram_reg_190__14_ ( .D(n7491), .CLK(clk), .Q(ram[3054]) );
  DFFPOSX1 ram_reg_190__13_ ( .D(n7490), .CLK(clk), .Q(ram[3053]) );
  DFFPOSX1 ram_reg_190__12_ ( .D(n7489), .CLK(clk), .Q(ram[3052]) );
  DFFPOSX1 ram_reg_190__11_ ( .D(n7488), .CLK(clk), .Q(ram[3051]) );
  DFFPOSX1 ram_reg_190__10_ ( .D(n7487), .CLK(clk), .Q(ram[3050]) );
  DFFPOSX1 ram_reg_190__9_ ( .D(n7486), .CLK(clk), .Q(ram[3049]) );
  DFFPOSX1 ram_reg_190__8_ ( .D(n7485), .CLK(clk), .Q(ram[3048]) );
  DFFPOSX1 ram_reg_190__7_ ( .D(n7484), .CLK(clk), .Q(ram[3047]) );
  DFFPOSX1 ram_reg_190__6_ ( .D(n7483), .CLK(clk), .Q(ram[3046]) );
  DFFPOSX1 ram_reg_190__5_ ( .D(n7482), .CLK(clk), .Q(ram[3045]) );
  DFFPOSX1 ram_reg_190__4_ ( .D(n7481), .CLK(clk), .Q(ram[3044]) );
  DFFPOSX1 ram_reg_190__3_ ( .D(n7480), .CLK(clk), .Q(ram[3043]) );
  DFFPOSX1 ram_reg_190__2_ ( .D(n7479), .CLK(clk), .Q(ram[3042]) );
  DFFPOSX1 ram_reg_190__1_ ( .D(n7478), .CLK(clk), .Q(ram[3041]) );
  DFFPOSX1 ram_reg_190__0_ ( .D(n7477), .CLK(clk), .Q(ram[3040]) );
  DFFPOSX1 ram_reg_189__15_ ( .D(n7476), .CLK(clk), .Q(ram[3039]) );
  DFFPOSX1 ram_reg_189__14_ ( .D(n7475), .CLK(clk), .Q(ram[3038]) );
  DFFPOSX1 ram_reg_189__13_ ( .D(n7474), .CLK(clk), .Q(ram[3037]) );
  DFFPOSX1 ram_reg_189__12_ ( .D(n7473), .CLK(clk), .Q(ram[3036]) );
  DFFPOSX1 ram_reg_189__11_ ( .D(n7472), .CLK(clk), .Q(ram[3035]) );
  DFFPOSX1 ram_reg_189__10_ ( .D(n7471), .CLK(clk), .Q(ram[3034]) );
  DFFPOSX1 ram_reg_189__9_ ( .D(n7470), .CLK(clk), .Q(ram[3033]) );
  DFFPOSX1 ram_reg_189__8_ ( .D(n7469), .CLK(clk), .Q(ram[3032]) );
  DFFPOSX1 ram_reg_189__7_ ( .D(n7468), .CLK(clk), .Q(ram[3031]) );
  DFFPOSX1 ram_reg_189__6_ ( .D(n7467), .CLK(clk), .Q(ram[3030]) );
  DFFPOSX1 ram_reg_189__5_ ( .D(n7466), .CLK(clk), .Q(ram[3029]) );
  DFFPOSX1 ram_reg_189__4_ ( .D(n7465), .CLK(clk), .Q(ram[3028]) );
  DFFPOSX1 ram_reg_189__3_ ( .D(n7464), .CLK(clk), .Q(ram[3027]) );
  DFFPOSX1 ram_reg_189__2_ ( .D(n7463), .CLK(clk), .Q(ram[3026]) );
  DFFPOSX1 ram_reg_189__1_ ( .D(n7462), .CLK(clk), .Q(ram[3025]) );
  DFFPOSX1 ram_reg_189__0_ ( .D(n7461), .CLK(clk), .Q(ram[3024]) );
  DFFPOSX1 ram_reg_188__15_ ( .D(n7460), .CLK(clk), .Q(ram[3023]) );
  DFFPOSX1 ram_reg_188__14_ ( .D(n7459), .CLK(clk), .Q(ram[3022]) );
  DFFPOSX1 ram_reg_188__13_ ( .D(n7458), .CLK(clk), .Q(ram[3021]) );
  DFFPOSX1 ram_reg_188__12_ ( .D(n7457), .CLK(clk), .Q(ram[3020]) );
  DFFPOSX1 ram_reg_188__11_ ( .D(n7456), .CLK(clk), .Q(ram[3019]) );
  DFFPOSX1 ram_reg_188__10_ ( .D(n7455), .CLK(clk), .Q(ram[3018]) );
  DFFPOSX1 ram_reg_188__9_ ( .D(n7454), .CLK(clk), .Q(ram[3017]) );
  DFFPOSX1 ram_reg_188__8_ ( .D(n7453), .CLK(clk), .Q(ram[3016]) );
  DFFPOSX1 ram_reg_188__7_ ( .D(n7452), .CLK(clk), .Q(ram[3015]) );
  DFFPOSX1 ram_reg_188__6_ ( .D(n7451), .CLK(clk), .Q(ram[3014]) );
  DFFPOSX1 ram_reg_188__5_ ( .D(n7450), .CLK(clk), .Q(ram[3013]) );
  DFFPOSX1 ram_reg_188__4_ ( .D(n7449), .CLK(clk), .Q(ram[3012]) );
  DFFPOSX1 ram_reg_188__3_ ( .D(n7448), .CLK(clk), .Q(ram[3011]) );
  DFFPOSX1 ram_reg_188__2_ ( .D(n7447), .CLK(clk), .Q(ram[3010]) );
  DFFPOSX1 ram_reg_188__1_ ( .D(n7446), .CLK(clk), .Q(ram[3009]) );
  DFFPOSX1 ram_reg_188__0_ ( .D(n7445), .CLK(clk), .Q(ram[3008]) );
  DFFPOSX1 ram_reg_187__15_ ( .D(n7444), .CLK(clk), .Q(ram[3007]) );
  DFFPOSX1 ram_reg_187__14_ ( .D(n7443), .CLK(clk), .Q(ram[3006]) );
  DFFPOSX1 ram_reg_187__13_ ( .D(n7442), .CLK(clk), .Q(ram[3005]) );
  DFFPOSX1 ram_reg_187__12_ ( .D(n7441), .CLK(clk), .Q(ram[3004]) );
  DFFPOSX1 ram_reg_187__11_ ( .D(n7440), .CLK(clk), .Q(ram[3003]) );
  DFFPOSX1 ram_reg_187__10_ ( .D(n7439), .CLK(clk), .Q(ram[3002]) );
  DFFPOSX1 ram_reg_187__9_ ( .D(n7438), .CLK(clk), .Q(ram[3001]) );
  DFFPOSX1 ram_reg_187__8_ ( .D(n7437), .CLK(clk), .Q(ram[3000]) );
  DFFPOSX1 ram_reg_187__7_ ( .D(n7436), .CLK(clk), .Q(ram[2999]) );
  DFFPOSX1 ram_reg_187__6_ ( .D(n7435), .CLK(clk), .Q(ram[2998]) );
  DFFPOSX1 ram_reg_187__5_ ( .D(n7434), .CLK(clk), .Q(ram[2997]) );
  DFFPOSX1 ram_reg_187__4_ ( .D(n7433), .CLK(clk), .Q(ram[2996]) );
  DFFPOSX1 ram_reg_187__3_ ( .D(n7432), .CLK(clk), .Q(ram[2995]) );
  DFFPOSX1 ram_reg_187__2_ ( .D(n7431), .CLK(clk), .Q(ram[2994]) );
  DFFPOSX1 ram_reg_187__1_ ( .D(n7430), .CLK(clk), .Q(ram[2993]) );
  DFFPOSX1 ram_reg_187__0_ ( .D(n7429), .CLK(clk), .Q(ram[2992]) );
  DFFPOSX1 ram_reg_186__15_ ( .D(n7428), .CLK(clk), .Q(ram[2991]) );
  DFFPOSX1 ram_reg_186__14_ ( .D(n7427), .CLK(clk), .Q(ram[2990]) );
  DFFPOSX1 ram_reg_186__13_ ( .D(n7426), .CLK(clk), .Q(ram[2989]) );
  DFFPOSX1 ram_reg_186__12_ ( .D(n7425), .CLK(clk), .Q(ram[2988]) );
  DFFPOSX1 ram_reg_186__11_ ( .D(n7424), .CLK(clk), .Q(ram[2987]) );
  DFFPOSX1 ram_reg_186__10_ ( .D(n7423), .CLK(clk), .Q(ram[2986]) );
  DFFPOSX1 ram_reg_186__9_ ( .D(n7422), .CLK(clk), .Q(ram[2985]) );
  DFFPOSX1 ram_reg_186__8_ ( .D(n7421), .CLK(clk), .Q(ram[2984]) );
  DFFPOSX1 ram_reg_186__7_ ( .D(n7420), .CLK(clk), .Q(ram[2983]) );
  DFFPOSX1 ram_reg_186__6_ ( .D(n7419), .CLK(clk), .Q(ram[2982]) );
  DFFPOSX1 ram_reg_186__5_ ( .D(n7418), .CLK(clk), .Q(ram[2981]) );
  DFFPOSX1 ram_reg_186__4_ ( .D(n7417), .CLK(clk), .Q(ram[2980]) );
  DFFPOSX1 ram_reg_186__3_ ( .D(n7416), .CLK(clk), .Q(ram[2979]) );
  DFFPOSX1 ram_reg_186__2_ ( .D(n7415), .CLK(clk), .Q(ram[2978]) );
  DFFPOSX1 ram_reg_186__1_ ( .D(n7414), .CLK(clk), .Q(ram[2977]) );
  DFFPOSX1 ram_reg_186__0_ ( .D(n7413), .CLK(clk), .Q(ram[2976]) );
  DFFPOSX1 ram_reg_185__15_ ( .D(n7412), .CLK(clk), .Q(ram[2975]) );
  DFFPOSX1 ram_reg_185__14_ ( .D(n7411), .CLK(clk), .Q(ram[2974]) );
  DFFPOSX1 ram_reg_185__13_ ( .D(n7410), .CLK(clk), .Q(ram[2973]) );
  DFFPOSX1 ram_reg_185__12_ ( .D(n7409), .CLK(clk), .Q(ram[2972]) );
  DFFPOSX1 ram_reg_185__11_ ( .D(n7408), .CLK(clk), .Q(ram[2971]) );
  DFFPOSX1 ram_reg_185__10_ ( .D(n7407), .CLK(clk), .Q(ram[2970]) );
  DFFPOSX1 ram_reg_185__9_ ( .D(n7406), .CLK(clk), .Q(ram[2969]) );
  DFFPOSX1 ram_reg_185__8_ ( .D(n7405), .CLK(clk), .Q(ram[2968]) );
  DFFPOSX1 ram_reg_185__7_ ( .D(n7404), .CLK(clk), .Q(ram[2967]) );
  DFFPOSX1 ram_reg_185__6_ ( .D(n7403), .CLK(clk), .Q(ram[2966]) );
  DFFPOSX1 ram_reg_185__5_ ( .D(n7402), .CLK(clk), .Q(ram[2965]) );
  DFFPOSX1 ram_reg_185__4_ ( .D(n7401), .CLK(clk), .Q(ram[2964]) );
  DFFPOSX1 ram_reg_185__3_ ( .D(n7400), .CLK(clk), .Q(ram[2963]) );
  DFFPOSX1 ram_reg_185__2_ ( .D(n7399), .CLK(clk), .Q(ram[2962]) );
  DFFPOSX1 ram_reg_185__1_ ( .D(n7398), .CLK(clk), .Q(ram[2961]) );
  DFFPOSX1 ram_reg_185__0_ ( .D(n7397), .CLK(clk), .Q(ram[2960]) );
  DFFPOSX1 ram_reg_184__15_ ( .D(n7396), .CLK(clk), .Q(ram[2959]) );
  DFFPOSX1 ram_reg_184__14_ ( .D(n7395), .CLK(clk), .Q(ram[2958]) );
  DFFPOSX1 ram_reg_184__13_ ( .D(n7394), .CLK(clk), .Q(ram[2957]) );
  DFFPOSX1 ram_reg_184__12_ ( .D(n7393), .CLK(clk), .Q(ram[2956]) );
  DFFPOSX1 ram_reg_184__11_ ( .D(n7392), .CLK(clk), .Q(ram[2955]) );
  DFFPOSX1 ram_reg_184__10_ ( .D(n7391), .CLK(clk), .Q(ram[2954]) );
  DFFPOSX1 ram_reg_184__9_ ( .D(n7390), .CLK(clk), .Q(ram[2953]) );
  DFFPOSX1 ram_reg_184__8_ ( .D(n7389), .CLK(clk), .Q(ram[2952]) );
  DFFPOSX1 ram_reg_184__7_ ( .D(n7388), .CLK(clk), .Q(ram[2951]) );
  DFFPOSX1 ram_reg_184__6_ ( .D(n7387), .CLK(clk), .Q(ram[2950]) );
  DFFPOSX1 ram_reg_184__5_ ( .D(n7386), .CLK(clk), .Q(ram[2949]) );
  DFFPOSX1 ram_reg_184__4_ ( .D(n7385), .CLK(clk), .Q(ram[2948]) );
  DFFPOSX1 ram_reg_184__3_ ( .D(n7384), .CLK(clk), .Q(ram[2947]) );
  DFFPOSX1 ram_reg_184__2_ ( .D(n7383), .CLK(clk), .Q(ram[2946]) );
  DFFPOSX1 ram_reg_184__1_ ( .D(n7382), .CLK(clk), .Q(ram[2945]) );
  DFFPOSX1 ram_reg_184__0_ ( .D(n7381), .CLK(clk), .Q(ram[2944]) );
  DFFPOSX1 ram_reg_183__15_ ( .D(n7380), .CLK(clk), .Q(ram[2943]) );
  DFFPOSX1 ram_reg_183__14_ ( .D(n7379), .CLK(clk), .Q(ram[2942]) );
  DFFPOSX1 ram_reg_183__13_ ( .D(n7378), .CLK(clk), .Q(ram[2941]) );
  DFFPOSX1 ram_reg_183__12_ ( .D(n7377), .CLK(clk), .Q(ram[2940]) );
  DFFPOSX1 ram_reg_183__11_ ( .D(n7376), .CLK(clk), .Q(ram[2939]) );
  DFFPOSX1 ram_reg_183__10_ ( .D(n7375), .CLK(clk), .Q(ram[2938]) );
  DFFPOSX1 ram_reg_183__9_ ( .D(n7374), .CLK(clk), .Q(ram[2937]) );
  DFFPOSX1 ram_reg_183__8_ ( .D(n7373), .CLK(clk), .Q(ram[2936]) );
  DFFPOSX1 ram_reg_183__7_ ( .D(n7372), .CLK(clk), .Q(ram[2935]) );
  DFFPOSX1 ram_reg_183__6_ ( .D(n7371), .CLK(clk), .Q(ram[2934]) );
  DFFPOSX1 ram_reg_183__5_ ( .D(n7370), .CLK(clk), .Q(ram[2933]) );
  DFFPOSX1 ram_reg_183__4_ ( .D(n7369), .CLK(clk), .Q(ram[2932]) );
  DFFPOSX1 ram_reg_183__3_ ( .D(n7368), .CLK(clk), .Q(ram[2931]) );
  DFFPOSX1 ram_reg_183__2_ ( .D(n7367), .CLK(clk), .Q(ram[2930]) );
  DFFPOSX1 ram_reg_183__1_ ( .D(n7366), .CLK(clk), .Q(ram[2929]) );
  DFFPOSX1 ram_reg_183__0_ ( .D(n7365), .CLK(clk), .Q(ram[2928]) );
  DFFPOSX1 ram_reg_182__15_ ( .D(n7364), .CLK(clk), .Q(ram[2927]) );
  DFFPOSX1 ram_reg_182__14_ ( .D(n7363), .CLK(clk), .Q(ram[2926]) );
  DFFPOSX1 ram_reg_182__13_ ( .D(n7362), .CLK(clk), .Q(ram[2925]) );
  DFFPOSX1 ram_reg_182__12_ ( .D(n7361), .CLK(clk), .Q(ram[2924]) );
  DFFPOSX1 ram_reg_182__11_ ( .D(n7360), .CLK(clk), .Q(ram[2923]) );
  DFFPOSX1 ram_reg_182__10_ ( .D(n7359), .CLK(clk), .Q(ram[2922]) );
  DFFPOSX1 ram_reg_182__9_ ( .D(n7358), .CLK(clk), .Q(ram[2921]) );
  DFFPOSX1 ram_reg_182__8_ ( .D(n7357), .CLK(clk), .Q(ram[2920]) );
  DFFPOSX1 ram_reg_182__7_ ( .D(n7356), .CLK(clk), .Q(ram[2919]) );
  DFFPOSX1 ram_reg_182__6_ ( .D(n7355), .CLK(clk), .Q(ram[2918]) );
  DFFPOSX1 ram_reg_182__5_ ( .D(n7354), .CLK(clk), .Q(ram[2917]) );
  DFFPOSX1 ram_reg_182__4_ ( .D(n7353), .CLK(clk), .Q(ram[2916]) );
  DFFPOSX1 ram_reg_182__3_ ( .D(n7352), .CLK(clk), .Q(ram[2915]) );
  DFFPOSX1 ram_reg_182__2_ ( .D(n7351), .CLK(clk), .Q(ram[2914]) );
  DFFPOSX1 ram_reg_182__1_ ( .D(n7350), .CLK(clk), .Q(ram[2913]) );
  DFFPOSX1 ram_reg_182__0_ ( .D(n7349), .CLK(clk), .Q(ram[2912]) );
  DFFPOSX1 ram_reg_181__15_ ( .D(n7348), .CLK(clk), .Q(ram[2911]) );
  DFFPOSX1 ram_reg_181__14_ ( .D(n7347), .CLK(clk), .Q(ram[2910]) );
  DFFPOSX1 ram_reg_181__13_ ( .D(n7346), .CLK(clk), .Q(ram[2909]) );
  DFFPOSX1 ram_reg_181__12_ ( .D(n7345), .CLK(clk), .Q(ram[2908]) );
  DFFPOSX1 ram_reg_181__11_ ( .D(n7344), .CLK(clk), .Q(ram[2907]) );
  DFFPOSX1 ram_reg_181__10_ ( .D(n7343), .CLK(clk), .Q(ram[2906]) );
  DFFPOSX1 ram_reg_181__9_ ( .D(n7342), .CLK(clk), .Q(ram[2905]) );
  DFFPOSX1 ram_reg_181__8_ ( .D(n7341), .CLK(clk), .Q(ram[2904]) );
  DFFPOSX1 ram_reg_181__7_ ( .D(n7340), .CLK(clk), .Q(ram[2903]) );
  DFFPOSX1 ram_reg_181__6_ ( .D(n7339), .CLK(clk), .Q(ram[2902]) );
  DFFPOSX1 ram_reg_181__5_ ( .D(n7338), .CLK(clk), .Q(ram[2901]) );
  DFFPOSX1 ram_reg_181__4_ ( .D(n7337), .CLK(clk), .Q(ram[2900]) );
  DFFPOSX1 ram_reg_181__3_ ( .D(n7336), .CLK(clk), .Q(ram[2899]) );
  DFFPOSX1 ram_reg_181__2_ ( .D(n7335), .CLK(clk), .Q(ram[2898]) );
  DFFPOSX1 ram_reg_181__1_ ( .D(n7334), .CLK(clk), .Q(ram[2897]) );
  DFFPOSX1 ram_reg_181__0_ ( .D(n7333), .CLK(clk), .Q(ram[2896]) );
  DFFPOSX1 ram_reg_180__15_ ( .D(n7332), .CLK(clk), .Q(ram[2895]) );
  DFFPOSX1 ram_reg_180__14_ ( .D(n7331), .CLK(clk), .Q(ram[2894]) );
  DFFPOSX1 ram_reg_180__13_ ( .D(n7330), .CLK(clk), .Q(ram[2893]) );
  DFFPOSX1 ram_reg_180__12_ ( .D(n7329), .CLK(clk), .Q(ram[2892]) );
  DFFPOSX1 ram_reg_180__11_ ( .D(n7328), .CLK(clk), .Q(ram[2891]) );
  DFFPOSX1 ram_reg_180__10_ ( .D(n7327), .CLK(clk), .Q(ram[2890]) );
  DFFPOSX1 ram_reg_180__9_ ( .D(n7326), .CLK(clk), .Q(ram[2889]) );
  DFFPOSX1 ram_reg_180__8_ ( .D(n7325), .CLK(clk), .Q(ram[2888]) );
  DFFPOSX1 ram_reg_180__7_ ( .D(n7324), .CLK(clk), .Q(ram[2887]) );
  DFFPOSX1 ram_reg_180__6_ ( .D(n7323), .CLK(clk), .Q(ram[2886]) );
  DFFPOSX1 ram_reg_180__5_ ( .D(n7322), .CLK(clk), .Q(ram[2885]) );
  DFFPOSX1 ram_reg_180__4_ ( .D(n7321), .CLK(clk), .Q(ram[2884]) );
  DFFPOSX1 ram_reg_180__3_ ( .D(n7320), .CLK(clk), .Q(ram[2883]) );
  DFFPOSX1 ram_reg_180__2_ ( .D(n7319), .CLK(clk), .Q(ram[2882]) );
  DFFPOSX1 ram_reg_180__1_ ( .D(n7318), .CLK(clk), .Q(ram[2881]) );
  DFFPOSX1 ram_reg_180__0_ ( .D(n7317), .CLK(clk), .Q(ram[2880]) );
  DFFPOSX1 ram_reg_179__15_ ( .D(n7316), .CLK(clk), .Q(ram[2879]) );
  DFFPOSX1 ram_reg_179__14_ ( .D(n7315), .CLK(clk), .Q(ram[2878]) );
  DFFPOSX1 ram_reg_179__13_ ( .D(n7314), .CLK(clk), .Q(ram[2877]) );
  DFFPOSX1 ram_reg_179__12_ ( .D(n7313), .CLK(clk), .Q(ram[2876]) );
  DFFPOSX1 ram_reg_179__11_ ( .D(n7312), .CLK(clk), .Q(ram[2875]) );
  DFFPOSX1 ram_reg_179__10_ ( .D(n7311), .CLK(clk), .Q(ram[2874]) );
  DFFPOSX1 ram_reg_179__9_ ( .D(n7310), .CLK(clk), .Q(ram[2873]) );
  DFFPOSX1 ram_reg_179__8_ ( .D(n7309), .CLK(clk), .Q(ram[2872]) );
  DFFPOSX1 ram_reg_179__7_ ( .D(n7308), .CLK(clk), .Q(ram[2871]) );
  DFFPOSX1 ram_reg_179__6_ ( .D(n7307), .CLK(clk), .Q(ram[2870]) );
  DFFPOSX1 ram_reg_179__5_ ( .D(n7306), .CLK(clk), .Q(ram[2869]) );
  DFFPOSX1 ram_reg_179__4_ ( .D(n7305), .CLK(clk), .Q(ram[2868]) );
  DFFPOSX1 ram_reg_179__3_ ( .D(n7304), .CLK(clk), .Q(ram[2867]) );
  DFFPOSX1 ram_reg_179__2_ ( .D(n7303), .CLK(clk), .Q(ram[2866]) );
  DFFPOSX1 ram_reg_179__1_ ( .D(n7302), .CLK(clk), .Q(ram[2865]) );
  DFFPOSX1 ram_reg_179__0_ ( .D(n7301), .CLK(clk), .Q(ram[2864]) );
  DFFPOSX1 ram_reg_178__15_ ( .D(n7300), .CLK(clk), .Q(ram[2863]) );
  DFFPOSX1 ram_reg_178__14_ ( .D(n7299), .CLK(clk), .Q(ram[2862]) );
  DFFPOSX1 ram_reg_178__13_ ( .D(n7298), .CLK(clk), .Q(ram[2861]) );
  DFFPOSX1 ram_reg_178__12_ ( .D(n7297), .CLK(clk), .Q(ram[2860]) );
  DFFPOSX1 ram_reg_178__11_ ( .D(n7296), .CLK(clk), .Q(ram[2859]) );
  DFFPOSX1 ram_reg_178__10_ ( .D(n7295), .CLK(clk), .Q(ram[2858]) );
  DFFPOSX1 ram_reg_178__9_ ( .D(n7294), .CLK(clk), .Q(ram[2857]) );
  DFFPOSX1 ram_reg_178__8_ ( .D(n7293), .CLK(clk), .Q(ram[2856]) );
  DFFPOSX1 ram_reg_178__7_ ( .D(n7292), .CLK(clk), .Q(ram[2855]) );
  DFFPOSX1 ram_reg_178__6_ ( .D(n7291), .CLK(clk), .Q(ram[2854]) );
  DFFPOSX1 ram_reg_178__5_ ( .D(n7290), .CLK(clk), .Q(ram[2853]) );
  DFFPOSX1 ram_reg_178__4_ ( .D(n7289), .CLK(clk), .Q(ram[2852]) );
  DFFPOSX1 ram_reg_178__3_ ( .D(n7288), .CLK(clk), .Q(ram[2851]) );
  DFFPOSX1 ram_reg_178__2_ ( .D(n7287), .CLK(clk), .Q(ram[2850]) );
  DFFPOSX1 ram_reg_178__1_ ( .D(n7286), .CLK(clk), .Q(ram[2849]) );
  DFFPOSX1 ram_reg_178__0_ ( .D(n7285), .CLK(clk), .Q(ram[2848]) );
  DFFPOSX1 ram_reg_177__15_ ( .D(n7284), .CLK(clk), .Q(ram[2847]) );
  DFFPOSX1 ram_reg_177__14_ ( .D(n7283), .CLK(clk), .Q(ram[2846]) );
  DFFPOSX1 ram_reg_177__13_ ( .D(n7282), .CLK(clk), .Q(ram[2845]) );
  DFFPOSX1 ram_reg_177__12_ ( .D(n7281), .CLK(clk), .Q(ram[2844]) );
  DFFPOSX1 ram_reg_177__11_ ( .D(n7280), .CLK(clk), .Q(ram[2843]) );
  DFFPOSX1 ram_reg_177__10_ ( .D(n7279), .CLK(clk), .Q(ram[2842]) );
  DFFPOSX1 ram_reg_177__9_ ( .D(n7278), .CLK(clk), .Q(ram[2841]) );
  DFFPOSX1 ram_reg_177__8_ ( .D(n7277), .CLK(clk), .Q(ram[2840]) );
  DFFPOSX1 ram_reg_177__7_ ( .D(n7276), .CLK(clk), .Q(ram[2839]) );
  DFFPOSX1 ram_reg_177__6_ ( .D(n7275), .CLK(clk), .Q(ram[2838]) );
  DFFPOSX1 ram_reg_177__5_ ( .D(n7274), .CLK(clk), .Q(ram[2837]) );
  DFFPOSX1 ram_reg_177__4_ ( .D(n7273), .CLK(clk), .Q(ram[2836]) );
  DFFPOSX1 ram_reg_177__3_ ( .D(n7272), .CLK(clk), .Q(ram[2835]) );
  DFFPOSX1 ram_reg_177__2_ ( .D(n7271), .CLK(clk), .Q(ram[2834]) );
  DFFPOSX1 ram_reg_177__1_ ( .D(n7270), .CLK(clk), .Q(ram[2833]) );
  DFFPOSX1 ram_reg_177__0_ ( .D(n7269), .CLK(clk), .Q(ram[2832]) );
  DFFPOSX1 ram_reg_176__15_ ( .D(n7268), .CLK(clk), .Q(ram[2831]) );
  DFFPOSX1 ram_reg_176__14_ ( .D(n7267), .CLK(clk), .Q(ram[2830]) );
  DFFPOSX1 ram_reg_176__13_ ( .D(n7266), .CLK(clk), .Q(ram[2829]) );
  DFFPOSX1 ram_reg_176__12_ ( .D(n7265), .CLK(clk), .Q(ram[2828]) );
  DFFPOSX1 ram_reg_176__11_ ( .D(n7264), .CLK(clk), .Q(ram[2827]) );
  DFFPOSX1 ram_reg_176__10_ ( .D(n7263), .CLK(clk), .Q(ram[2826]) );
  DFFPOSX1 ram_reg_176__9_ ( .D(n7262), .CLK(clk), .Q(ram[2825]) );
  DFFPOSX1 ram_reg_176__8_ ( .D(n7261), .CLK(clk), .Q(ram[2824]) );
  DFFPOSX1 ram_reg_176__7_ ( .D(n7260), .CLK(clk), .Q(ram[2823]) );
  DFFPOSX1 ram_reg_176__6_ ( .D(n7259), .CLK(clk), .Q(ram[2822]) );
  DFFPOSX1 ram_reg_176__5_ ( .D(n7258), .CLK(clk), .Q(ram[2821]) );
  DFFPOSX1 ram_reg_176__4_ ( .D(n7257), .CLK(clk), .Q(ram[2820]) );
  DFFPOSX1 ram_reg_176__3_ ( .D(n7256), .CLK(clk), .Q(ram[2819]) );
  DFFPOSX1 ram_reg_176__2_ ( .D(n7255), .CLK(clk), .Q(ram[2818]) );
  DFFPOSX1 ram_reg_176__1_ ( .D(n7254), .CLK(clk), .Q(ram[2817]) );
  DFFPOSX1 ram_reg_176__0_ ( .D(n7253), .CLK(clk), .Q(ram[2816]) );
  DFFPOSX1 ram_reg_175__15_ ( .D(n7252), .CLK(clk), .Q(ram[2815]) );
  DFFPOSX1 ram_reg_175__14_ ( .D(n7251), .CLK(clk), .Q(ram[2814]) );
  DFFPOSX1 ram_reg_175__13_ ( .D(n7250), .CLK(clk), .Q(ram[2813]) );
  DFFPOSX1 ram_reg_175__12_ ( .D(n7249), .CLK(clk), .Q(ram[2812]) );
  DFFPOSX1 ram_reg_175__11_ ( .D(n7248), .CLK(clk), .Q(ram[2811]) );
  DFFPOSX1 ram_reg_175__10_ ( .D(n7247), .CLK(clk), .Q(ram[2810]) );
  DFFPOSX1 ram_reg_175__9_ ( .D(n7246), .CLK(clk), .Q(ram[2809]) );
  DFFPOSX1 ram_reg_175__8_ ( .D(n7245), .CLK(clk), .Q(ram[2808]) );
  DFFPOSX1 ram_reg_175__7_ ( .D(n7244), .CLK(clk), .Q(ram[2807]) );
  DFFPOSX1 ram_reg_175__6_ ( .D(n7243), .CLK(clk), .Q(ram[2806]) );
  DFFPOSX1 ram_reg_175__5_ ( .D(n7242), .CLK(clk), .Q(ram[2805]) );
  DFFPOSX1 ram_reg_175__4_ ( .D(n7241), .CLK(clk), .Q(ram[2804]) );
  DFFPOSX1 ram_reg_175__3_ ( .D(n7240), .CLK(clk), .Q(ram[2803]) );
  DFFPOSX1 ram_reg_175__2_ ( .D(n7239), .CLK(clk), .Q(ram[2802]) );
  DFFPOSX1 ram_reg_175__1_ ( .D(n7238), .CLK(clk), .Q(ram[2801]) );
  DFFPOSX1 ram_reg_175__0_ ( .D(n7237), .CLK(clk), .Q(ram[2800]) );
  DFFPOSX1 ram_reg_174__15_ ( .D(n7236), .CLK(clk), .Q(ram[2799]) );
  DFFPOSX1 ram_reg_174__14_ ( .D(n7235), .CLK(clk), .Q(ram[2798]) );
  DFFPOSX1 ram_reg_174__13_ ( .D(n7234), .CLK(clk), .Q(ram[2797]) );
  DFFPOSX1 ram_reg_174__12_ ( .D(n7233), .CLK(clk), .Q(ram[2796]) );
  DFFPOSX1 ram_reg_174__11_ ( .D(n7232), .CLK(clk), .Q(ram[2795]) );
  DFFPOSX1 ram_reg_174__10_ ( .D(n7231), .CLK(clk), .Q(ram[2794]) );
  DFFPOSX1 ram_reg_174__9_ ( .D(n7230), .CLK(clk), .Q(ram[2793]) );
  DFFPOSX1 ram_reg_174__8_ ( .D(n7229), .CLK(clk), .Q(ram[2792]) );
  DFFPOSX1 ram_reg_174__7_ ( .D(n7228), .CLK(clk), .Q(ram[2791]) );
  DFFPOSX1 ram_reg_174__6_ ( .D(n7227), .CLK(clk), .Q(ram[2790]) );
  DFFPOSX1 ram_reg_174__5_ ( .D(n7226), .CLK(clk), .Q(ram[2789]) );
  DFFPOSX1 ram_reg_174__4_ ( .D(n7225), .CLK(clk), .Q(ram[2788]) );
  DFFPOSX1 ram_reg_174__3_ ( .D(n7224), .CLK(clk), .Q(ram[2787]) );
  DFFPOSX1 ram_reg_174__2_ ( .D(n7223), .CLK(clk), .Q(ram[2786]) );
  DFFPOSX1 ram_reg_174__1_ ( .D(n7222), .CLK(clk), .Q(ram[2785]) );
  DFFPOSX1 ram_reg_174__0_ ( .D(n7221), .CLK(clk), .Q(ram[2784]) );
  DFFPOSX1 ram_reg_173__15_ ( .D(n7220), .CLK(clk), .Q(ram[2783]) );
  DFFPOSX1 ram_reg_173__14_ ( .D(n7219), .CLK(clk), .Q(ram[2782]) );
  DFFPOSX1 ram_reg_173__13_ ( .D(n7218), .CLK(clk), .Q(ram[2781]) );
  DFFPOSX1 ram_reg_173__12_ ( .D(n7217), .CLK(clk), .Q(ram[2780]) );
  DFFPOSX1 ram_reg_173__11_ ( .D(n7216), .CLK(clk), .Q(ram[2779]) );
  DFFPOSX1 ram_reg_173__10_ ( .D(n7215), .CLK(clk), .Q(ram[2778]) );
  DFFPOSX1 ram_reg_173__9_ ( .D(n7214), .CLK(clk), .Q(ram[2777]) );
  DFFPOSX1 ram_reg_173__8_ ( .D(n7213), .CLK(clk), .Q(ram[2776]) );
  DFFPOSX1 ram_reg_173__7_ ( .D(n7212), .CLK(clk), .Q(ram[2775]) );
  DFFPOSX1 ram_reg_173__6_ ( .D(n7211), .CLK(clk), .Q(ram[2774]) );
  DFFPOSX1 ram_reg_173__5_ ( .D(n7210), .CLK(clk), .Q(ram[2773]) );
  DFFPOSX1 ram_reg_173__4_ ( .D(n7209), .CLK(clk), .Q(ram[2772]) );
  DFFPOSX1 ram_reg_173__3_ ( .D(n7208), .CLK(clk), .Q(ram[2771]) );
  DFFPOSX1 ram_reg_173__2_ ( .D(n7207), .CLK(clk), .Q(ram[2770]) );
  DFFPOSX1 ram_reg_173__1_ ( .D(n7206), .CLK(clk), .Q(ram[2769]) );
  DFFPOSX1 ram_reg_173__0_ ( .D(n7205), .CLK(clk), .Q(ram[2768]) );
  DFFPOSX1 ram_reg_172__15_ ( .D(n7204), .CLK(clk), .Q(ram[2767]) );
  DFFPOSX1 ram_reg_172__14_ ( .D(n7203), .CLK(clk), .Q(ram[2766]) );
  DFFPOSX1 ram_reg_172__13_ ( .D(n7202), .CLK(clk), .Q(ram[2765]) );
  DFFPOSX1 ram_reg_172__12_ ( .D(n7201), .CLK(clk), .Q(ram[2764]) );
  DFFPOSX1 ram_reg_172__11_ ( .D(n7200), .CLK(clk), .Q(ram[2763]) );
  DFFPOSX1 ram_reg_172__10_ ( .D(n7199), .CLK(clk), .Q(ram[2762]) );
  DFFPOSX1 ram_reg_172__9_ ( .D(n7198), .CLK(clk), .Q(ram[2761]) );
  DFFPOSX1 ram_reg_172__8_ ( .D(n7197), .CLK(clk), .Q(ram[2760]) );
  DFFPOSX1 ram_reg_172__7_ ( .D(n7196), .CLK(clk), .Q(ram[2759]) );
  DFFPOSX1 ram_reg_172__6_ ( .D(n7195), .CLK(clk), .Q(ram[2758]) );
  DFFPOSX1 ram_reg_172__5_ ( .D(n7194), .CLK(clk), .Q(ram[2757]) );
  DFFPOSX1 ram_reg_172__4_ ( .D(n7193), .CLK(clk), .Q(ram[2756]) );
  DFFPOSX1 ram_reg_172__3_ ( .D(n7192), .CLK(clk), .Q(ram[2755]) );
  DFFPOSX1 ram_reg_172__2_ ( .D(n7191), .CLK(clk), .Q(ram[2754]) );
  DFFPOSX1 ram_reg_172__1_ ( .D(n7190), .CLK(clk), .Q(ram[2753]) );
  DFFPOSX1 ram_reg_172__0_ ( .D(n7189), .CLK(clk), .Q(ram[2752]) );
  DFFPOSX1 ram_reg_171__15_ ( .D(n7188), .CLK(clk), .Q(ram[2751]) );
  DFFPOSX1 ram_reg_171__14_ ( .D(n7187), .CLK(clk), .Q(ram[2750]) );
  DFFPOSX1 ram_reg_171__13_ ( .D(n7186), .CLK(clk), .Q(ram[2749]) );
  DFFPOSX1 ram_reg_171__12_ ( .D(n7185), .CLK(clk), .Q(ram[2748]) );
  DFFPOSX1 ram_reg_171__11_ ( .D(n7184), .CLK(clk), .Q(ram[2747]) );
  DFFPOSX1 ram_reg_171__10_ ( .D(n7183), .CLK(clk), .Q(ram[2746]) );
  DFFPOSX1 ram_reg_171__9_ ( .D(n7182), .CLK(clk), .Q(ram[2745]) );
  DFFPOSX1 ram_reg_171__8_ ( .D(n7181), .CLK(clk), .Q(ram[2744]) );
  DFFPOSX1 ram_reg_171__7_ ( .D(n7180), .CLK(clk), .Q(ram[2743]) );
  DFFPOSX1 ram_reg_171__6_ ( .D(n7179), .CLK(clk), .Q(ram[2742]) );
  DFFPOSX1 ram_reg_171__5_ ( .D(n7178), .CLK(clk), .Q(ram[2741]) );
  DFFPOSX1 ram_reg_171__4_ ( .D(n7177), .CLK(clk), .Q(ram[2740]) );
  DFFPOSX1 ram_reg_171__3_ ( .D(n7176), .CLK(clk), .Q(ram[2739]) );
  DFFPOSX1 ram_reg_171__2_ ( .D(n7175), .CLK(clk), .Q(ram[2738]) );
  DFFPOSX1 ram_reg_171__1_ ( .D(n7174), .CLK(clk), .Q(ram[2737]) );
  DFFPOSX1 ram_reg_171__0_ ( .D(n7173), .CLK(clk), .Q(ram[2736]) );
  DFFPOSX1 ram_reg_170__15_ ( .D(n7172), .CLK(clk), .Q(ram[2735]) );
  DFFPOSX1 ram_reg_170__14_ ( .D(n7171), .CLK(clk), .Q(ram[2734]) );
  DFFPOSX1 ram_reg_170__13_ ( .D(n7170), .CLK(clk), .Q(ram[2733]) );
  DFFPOSX1 ram_reg_170__12_ ( .D(n7169), .CLK(clk), .Q(ram[2732]) );
  DFFPOSX1 ram_reg_170__11_ ( .D(n7168), .CLK(clk), .Q(ram[2731]) );
  DFFPOSX1 ram_reg_170__10_ ( .D(n7167), .CLK(clk), .Q(ram[2730]) );
  DFFPOSX1 ram_reg_170__9_ ( .D(n7166), .CLK(clk), .Q(ram[2729]) );
  DFFPOSX1 ram_reg_170__8_ ( .D(n7165), .CLK(clk), .Q(ram[2728]) );
  DFFPOSX1 ram_reg_170__7_ ( .D(n7164), .CLK(clk), .Q(ram[2727]) );
  DFFPOSX1 ram_reg_170__6_ ( .D(n7163), .CLK(clk), .Q(ram[2726]) );
  DFFPOSX1 ram_reg_170__5_ ( .D(n7162), .CLK(clk), .Q(ram[2725]) );
  DFFPOSX1 ram_reg_170__4_ ( .D(n7161), .CLK(clk), .Q(ram[2724]) );
  DFFPOSX1 ram_reg_170__3_ ( .D(n7160), .CLK(clk), .Q(ram[2723]) );
  DFFPOSX1 ram_reg_170__2_ ( .D(n7159), .CLK(clk), .Q(ram[2722]) );
  DFFPOSX1 ram_reg_170__1_ ( .D(n7158), .CLK(clk), .Q(ram[2721]) );
  DFFPOSX1 ram_reg_170__0_ ( .D(n7157), .CLK(clk), .Q(ram[2720]) );
  DFFPOSX1 ram_reg_169__15_ ( .D(n7156), .CLK(clk), .Q(ram[2719]) );
  DFFPOSX1 ram_reg_169__14_ ( .D(n7155), .CLK(clk), .Q(ram[2718]) );
  DFFPOSX1 ram_reg_169__13_ ( .D(n7154), .CLK(clk), .Q(ram[2717]) );
  DFFPOSX1 ram_reg_169__12_ ( .D(n7153), .CLK(clk), .Q(ram[2716]) );
  DFFPOSX1 ram_reg_169__11_ ( .D(n7152), .CLK(clk), .Q(ram[2715]) );
  DFFPOSX1 ram_reg_169__10_ ( .D(n7151), .CLK(clk), .Q(ram[2714]) );
  DFFPOSX1 ram_reg_169__9_ ( .D(n7150), .CLK(clk), .Q(ram[2713]) );
  DFFPOSX1 ram_reg_169__8_ ( .D(n7149), .CLK(clk), .Q(ram[2712]) );
  DFFPOSX1 ram_reg_169__7_ ( .D(n7148), .CLK(clk), .Q(ram[2711]) );
  DFFPOSX1 ram_reg_169__6_ ( .D(n7147), .CLK(clk), .Q(ram[2710]) );
  DFFPOSX1 ram_reg_169__5_ ( .D(n7146), .CLK(clk), .Q(ram[2709]) );
  DFFPOSX1 ram_reg_169__4_ ( .D(n7145), .CLK(clk), .Q(ram[2708]) );
  DFFPOSX1 ram_reg_169__3_ ( .D(n7144), .CLK(clk), .Q(ram[2707]) );
  DFFPOSX1 ram_reg_169__2_ ( .D(n7143), .CLK(clk), .Q(ram[2706]) );
  DFFPOSX1 ram_reg_169__1_ ( .D(n7142), .CLK(clk), .Q(ram[2705]) );
  DFFPOSX1 ram_reg_169__0_ ( .D(n7141), .CLK(clk), .Q(ram[2704]) );
  DFFPOSX1 ram_reg_168__15_ ( .D(n7140), .CLK(clk), .Q(ram[2703]) );
  DFFPOSX1 ram_reg_168__14_ ( .D(n7139), .CLK(clk), .Q(ram[2702]) );
  DFFPOSX1 ram_reg_168__13_ ( .D(n7138), .CLK(clk), .Q(ram[2701]) );
  DFFPOSX1 ram_reg_168__12_ ( .D(n7137), .CLK(clk), .Q(ram[2700]) );
  DFFPOSX1 ram_reg_168__11_ ( .D(n7136), .CLK(clk), .Q(ram[2699]) );
  DFFPOSX1 ram_reg_168__10_ ( .D(n7135), .CLK(clk), .Q(ram[2698]) );
  DFFPOSX1 ram_reg_168__9_ ( .D(n7134), .CLK(clk), .Q(ram[2697]) );
  DFFPOSX1 ram_reg_168__8_ ( .D(n7133), .CLK(clk), .Q(ram[2696]) );
  DFFPOSX1 ram_reg_168__7_ ( .D(n7132), .CLK(clk), .Q(ram[2695]) );
  DFFPOSX1 ram_reg_168__6_ ( .D(n7131), .CLK(clk), .Q(ram[2694]) );
  DFFPOSX1 ram_reg_168__5_ ( .D(n7130), .CLK(clk), .Q(ram[2693]) );
  DFFPOSX1 ram_reg_168__4_ ( .D(n7129), .CLK(clk), .Q(ram[2692]) );
  DFFPOSX1 ram_reg_168__3_ ( .D(n7128), .CLK(clk), .Q(ram[2691]) );
  DFFPOSX1 ram_reg_168__2_ ( .D(n7127), .CLK(clk), .Q(ram[2690]) );
  DFFPOSX1 ram_reg_168__1_ ( .D(n7126), .CLK(clk), .Q(ram[2689]) );
  DFFPOSX1 ram_reg_168__0_ ( .D(n7125), .CLK(clk), .Q(ram[2688]) );
  DFFPOSX1 ram_reg_167__15_ ( .D(n7124), .CLK(clk), .Q(ram[2687]) );
  DFFPOSX1 ram_reg_167__14_ ( .D(n7123), .CLK(clk), .Q(ram[2686]) );
  DFFPOSX1 ram_reg_167__13_ ( .D(n7122), .CLK(clk), .Q(ram[2685]) );
  DFFPOSX1 ram_reg_167__12_ ( .D(n7121), .CLK(clk), .Q(ram[2684]) );
  DFFPOSX1 ram_reg_167__11_ ( .D(n7120), .CLK(clk), .Q(ram[2683]) );
  DFFPOSX1 ram_reg_167__10_ ( .D(n7119), .CLK(clk), .Q(ram[2682]) );
  DFFPOSX1 ram_reg_167__9_ ( .D(n7118), .CLK(clk), .Q(ram[2681]) );
  DFFPOSX1 ram_reg_167__8_ ( .D(n7117), .CLK(clk), .Q(ram[2680]) );
  DFFPOSX1 ram_reg_167__7_ ( .D(n7116), .CLK(clk), .Q(ram[2679]) );
  DFFPOSX1 ram_reg_167__6_ ( .D(n7115), .CLK(clk), .Q(ram[2678]) );
  DFFPOSX1 ram_reg_167__5_ ( .D(n7114), .CLK(clk), .Q(ram[2677]) );
  DFFPOSX1 ram_reg_167__4_ ( .D(n7113), .CLK(clk), .Q(ram[2676]) );
  DFFPOSX1 ram_reg_167__3_ ( .D(n7112), .CLK(clk), .Q(ram[2675]) );
  DFFPOSX1 ram_reg_167__2_ ( .D(n7111), .CLK(clk), .Q(ram[2674]) );
  DFFPOSX1 ram_reg_167__1_ ( .D(n7110), .CLK(clk), .Q(ram[2673]) );
  DFFPOSX1 ram_reg_167__0_ ( .D(n7109), .CLK(clk), .Q(ram[2672]) );
  DFFPOSX1 ram_reg_166__15_ ( .D(n7108), .CLK(clk), .Q(ram[2671]) );
  DFFPOSX1 ram_reg_166__14_ ( .D(n7107), .CLK(clk), .Q(ram[2670]) );
  DFFPOSX1 ram_reg_166__13_ ( .D(n7106), .CLK(clk), .Q(ram[2669]) );
  DFFPOSX1 ram_reg_166__12_ ( .D(n7105), .CLK(clk), .Q(ram[2668]) );
  DFFPOSX1 ram_reg_166__11_ ( .D(n7104), .CLK(clk), .Q(ram[2667]) );
  DFFPOSX1 ram_reg_166__10_ ( .D(n7103), .CLK(clk), .Q(ram[2666]) );
  DFFPOSX1 ram_reg_166__9_ ( .D(n7102), .CLK(clk), .Q(ram[2665]) );
  DFFPOSX1 ram_reg_166__8_ ( .D(n7101), .CLK(clk), .Q(ram[2664]) );
  DFFPOSX1 ram_reg_166__7_ ( .D(n7100), .CLK(clk), .Q(ram[2663]) );
  DFFPOSX1 ram_reg_166__6_ ( .D(n7099), .CLK(clk), .Q(ram[2662]) );
  DFFPOSX1 ram_reg_166__5_ ( .D(n7098), .CLK(clk), .Q(ram[2661]) );
  DFFPOSX1 ram_reg_166__4_ ( .D(n7097), .CLK(clk), .Q(ram[2660]) );
  DFFPOSX1 ram_reg_166__3_ ( .D(n7096), .CLK(clk), .Q(ram[2659]) );
  DFFPOSX1 ram_reg_166__2_ ( .D(n7095), .CLK(clk), .Q(ram[2658]) );
  DFFPOSX1 ram_reg_166__1_ ( .D(n7094), .CLK(clk), .Q(ram[2657]) );
  DFFPOSX1 ram_reg_166__0_ ( .D(n7093), .CLK(clk), .Q(ram[2656]) );
  DFFPOSX1 ram_reg_165__15_ ( .D(n7092), .CLK(clk), .Q(ram[2655]) );
  DFFPOSX1 ram_reg_165__14_ ( .D(n7091), .CLK(clk), .Q(ram[2654]) );
  DFFPOSX1 ram_reg_165__13_ ( .D(n7090), .CLK(clk), .Q(ram[2653]) );
  DFFPOSX1 ram_reg_165__12_ ( .D(n7089), .CLK(clk), .Q(ram[2652]) );
  DFFPOSX1 ram_reg_165__11_ ( .D(n7088), .CLK(clk), .Q(ram[2651]) );
  DFFPOSX1 ram_reg_165__10_ ( .D(n7087), .CLK(clk), .Q(ram[2650]) );
  DFFPOSX1 ram_reg_165__9_ ( .D(n7086), .CLK(clk), .Q(ram[2649]) );
  DFFPOSX1 ram_reg_165__8_ ( .D(n7085), .CLK(clk), .Q(ram[2648]) );
  DFFPOSX1 ram_reg_165__7_ ( .D(n7084), .CLK(clk), .Q(ram[2647]) );
  DFFPOSX1 ram_reg_165__6_ ( .D(n7083), .CLK(clk), .Q(ram[2646]) );
  DFFPOSX1 ram_reg_165__5_ ( .D(n7082), .CLK(clk), .Q(ram[2645]) );
  DFFPOSX1 ram_reg_165__4_ ( .D(n7081), .CLK(clk), .Q(ram[2644]) );
  DFFPOSX1 ram_reg_165__3_ ( .D(n7080), .CLK(clk), .Q(ram[2643]) );
  DFFPOSX1 ram_reg_165__2_ ( .D(n7079), .CLK(clk), .Q(ram[2642]) );
  DFFPOSX1 ram_reg_165__1_ ( .D(n7078), .CLK(clk), .Q(ram[2641]) );
  DFFPOSX1 ram_reg_165__0_ ( .D(n7077), .CLK(clk), .Q(ram[2640]) );
  DFFPOSX1 ram_reg_164__15_ ( .D(n7076), .CLK(clk), .Q(ram[2639]) );
  DFFPOSX1 ram_reg_164__14_ ( .D(n7075), .CLK(clk), .Q(ram[2638]) );
  DFFPOSX1 ram_reg_164__13_ ( .D(n7074), .CLK(clk), .Q(ram[2637]) );
  DFFPOSX1 ram_reg_164__12_ ( .D(n7073), .CLK(clk), .Q(ram[2636]) );
  DFFPOSX1 ram_reg_164__11_ ( .D(n7072), .CLK(clk), .Q(ram[2635]) );
  DFFPOSX1 ram_reg_164__10_ ( .D(n7071), .CLK(clk), .Q(ram[2634]) );
  DFFPOSX1 ram_reg_164__9_ ( .D(n7070), .CLK(clk), .Q(ram[2633]) );
  DFFPOSX1 ram_reg_164__8_ ( .D(n7069), .CLK(clk), .Q(ram[2632]) );
  DFFPOSX1 ram_reg_164__7_ ( .D(n7068), .CLK(clk), .Q(ram[2631]) );
  DFFPOSX1 ram_reg_164__6_ ( .D(n7067), .CLK(clk), .Q(ram[2630]) );
  DFFPOSX1 ram_reg_164__5_ ( .D(n7066), .CLK(clk), .Q(ram[2629]) );
  DFFPOSX1 ram_reg_164__4_ ( .D(n7065), .CLK(clk), .Q(ram[2628]) );
  DFFPOSX1 ram_reg_164__3_ ( .D(n7064), .CLK(clk), .Q(ram[2627]) );
  DFFPOSX1 ram_reg_164__2_ ( .D(n7063), .CLK(clk), .Q(ram[2626]) );
  DFFPOSX1 ram_reg_164__1_ ( .D(n7062), .CLK(clk), .Q(ram[2625]) );
  DFFPOSX1 ram_reg_164__0_ ( .D(n7061), .CLK(clk), .Q(ram[2624]) );
  DFFPOSX1 ram_reg_163__15_ ( .D(n7060), .CLK(clk), .Q(ram[2623]) );
  DFFPOSX1 ram_reg_163__14_ ( .D(n7059), .CLK(clk), .Q(ram[2622]) );
  DFFPOSX1 ram_reg_163__13_ ( .D(n7058), .CLK(clk), .Q(ram[2621]) );
  DFFPOSX1 ram_reg_163__12_ ( .D(n7057), .CLK(clk), .Q(ram[2620]) );
  DFFPOSX1 ram_reg_163__11_ ( .D(n7056), .CLK(clk), .Q(ram[2619]) );
  DFFPOSX1 ram_reg_163__10_ ( .D(n7055), .CLK(clk), .Q(ram[2618]) );
  DFFPOSX1 ram_reg_163__9_ ( .D(n7054), .CLK(clk), .Q(ram[2617]) );
  DFFPOSX1 ram_reg_163__8_ ( .D(n7053), .CLK(clk), .Q(ram[2616]) );
  DFFPOSX1 ram_reg_163__7_ ( .D(n7052), .CLK(clk), .Q(ram[2615]) );
  DFFPOSX1 ram_reg_163__6_ ( .D(n7051), .CLK(clk), .Q(ram[2614]) );
  DFFPOSX1 ram_reg_163__5_ ( .D(n7050), .CLK(clk), .Q(ram[2613]) );
  DFFPOSX1 ram_reg_163__4_ ( .D(n7049), .CLK(clk), .Q(ram[2612]) );
  DFFPOSX1 ram_reg_163__3_ ( .D(n7048), .CLK(clk), .Q(ram[2611]) );
  DFFPOSX1 ram_reg_163__2_ ( .D(n7047), .CLK(clk), .Q(ram[2610]) );
  DFFPOSX1 ram_reg_163__1_ ( .D(n7046), .CLK(clk), .Q(ram[2609]) );
  DFFPOSX1 ram_reg_163__0_ ( .D(n7045), .CLK(clk), .Q(ram[2608]) );
  DFFPOSX1 ram_reg_162__15_ ( .D(n7044), .CLK(clk), .Q(ram[2607]) );
  DFFPOSX1 ram_reg_162__14_ ( .D(n7043), .CLK(clk), .Q(ram[2606]) );
  DFFPOSX1 ram_reg_162__13_ ( .D(n7042), .CLK(clk), .Q(ram[2605]) );
  DFFPOSX1 ram_reg_162__12_ ( .D(n7041), .CLK(clk), .Q(ram[2604]) );
  DFFPOSX1 ram_reg_162__11_ ( .D(n7040), .CLK(clk), .Q(ram[2603]) );
  DFFPOSX1 ram_reg_162__10_ ( .D(n7039), .CLK(clk), .Q(ram[2602]) );
  DFFPOSX1 ram_reg_162__9_ ( .D(n7038), .CLK(clk), .Q(ram[2601]) );
  DFFPOSX1 ram_reg_162__8_ ( .D(n7037), .CLK(clk), .Q(ram[2600]) );
  DFFPOSX1 ram_reg_162__7_ ( .D(n7036), .CLK(clk), .Q(ram[2599]) );
  DFFPOSX1 ram_reg_162__6_ ( .D(n7035), .CLK(clk), .Q(ram[2598]) );
  DFFPOSX1 ram_reg_162__5_ ( .D(n7034), .CLK(clk), .Q(ram[2597]) );
  DFFPOSX1 ram_reg_162__4_ ( .D(n7033), .CLK(clk), .Q(ram[2596]) );
  DFFPOSX1 ram_reg_162__3_ ( .D(n7032), .CLK(clk), .Q(ram[2595]) );
  DFFPOSX1 ram_reg_162__2_ ( .D(n7031), .CLK(clk), .Q(ram[2594]) );
  DFFPOSX1 ram_reg_162__1_ ( .D(n7030), .CLK(clk), .Q(ram[2593]) );
  DFFPOSX1 ram_reg_162__0_ ( .D(n7029), .CLK(clk), .Q(ram[2592]) );
  DFFPOSX1 ram_reg_161__15_ ( .D(n7028), .CLK(clk), .Q(ram[2591]) );
  DFFPOSX1 ram_reg_161__14_ ( .D(n7027), .CLK(clk), .Q(ram[2590]) );
  DFFPOSX1 ram_reg_161__13_ ( .D(n7026), .CLK(clk), .Q(ram[2589]) );
  DFFPOSX1 ram_reg_161__12_ ( .D(n7025), .CLK(clk), .Q(ram[2588]) );
  DFFPOSX1 ram_reg_161__11_ ( .D(n7024), .CLK(clk), .Q(ram[2587]) );
  DFFPOSX1 ram_reg_161__10_ ( .D(n7023), .CLK(clk), .Q(ram[2586]) );
  DFFPOSX1 ram_reg_161__9_ ( .D(n7022), .CLK(clk), .Q(ram[2585]) );
  DFFPOSX1 ram_reg_161__8_ ( .D(n7021), .CLK(clk), .Q(ram[2584]) );
  DFFPOSX1 ram_reg_161__7_ ( .D(n7020), .CLK(clk), .Q(ram[2583]) );
  DFFPOSX1 ram_reg_161__6_ ( .D(n7019), .CLK(clk), .Q(ram[2582]) );
  DFFPOSX1 ram_reg_161__5_ ( .D(n7018), .CLK(clk), .Q(ram[2581]) );
  DFFPOSX1 ram_reg_161__4_ ( .D(n7017), .CLK(clk), .Q(ram[2580]) );
  DFFPOSX1 ram_reg_161__3_ ( .D(n7016), .CLK(clk), .Q(ram[2579]) );
  DFFPOSX1 ram_reg_161__2_ ( .D(n7015), .CLK(clk), .Q(ram[2578]) );
  DFFPOSX1 ram_reg_161__1_ ( .D(n7014), .CLK(clk), .Q(ram[2577]) );
  DFFPOSX1 ram_reg_161__0_ ( .D(n7013), .CLK(clk), .Q(ram[2576]) );
  DFFPOSX1 ram_reg_160__15_ ( .D(n7012), .CLK(clk), .Q(ram[2575]) );
  DFFPOSX1 ram_reg_160__14_ ( .D(n7011), .CLK(clk), .Q(ram[2574]) );
  DFFPOSX1 ram_reg_160__13_ ( .D(n7010), .CLK(clk), .Q(ram[2573]) );
  DFFPOSX1 ram_reg_160__12_ ( .D(n7009), .CLK(clk), .Q(ram[2572]) );
  DFFPOSX1 ram_reg_160__11_ ( .D(n7008), .CLK(clk), .Q(ram[2571]) );
  DFFPOSX1 ram_reg_160__10_ ( .D(n7007), .CLK(clk), .Q(ram[2570]) );
  DFFPOSX1 ram_reg_160__9_ ( .D(n7006), .CLK(clk), .Q(ram[2569]) );
  DFFPOSX1 ram_reg_160__8_ ( .D(n7005), .CLK(clk), .Q(ram[2568]) );
  DFFPOSX1 ram_reg_160__7_ ( .D(n7004), .CLK(clk), .Q(ram[2567]) );
  DFFPOSX1 ram_reg_160__6_ ( .D(n7003), .CLK(clk), .Q(ram[2566]) );
  DFFPOSX1 ram_reg_160__5_ ( .D(n7002), .CLK(clk), .Q(ram[2565]) );
  DFFPOSX1 ram_reg_160__4_ ( .D(n7001), .CLK(clk), .Q(ram[2564]) );
  DFFPOSX1 ram_reg_160__3_ ( .D(n7000), .CLK(clk), .Q(ram[2563]) );
  DFFPOSX1 ram_reg_160__2_ ( .D(n6999), .CLK(clk), .Q(ram[2562]) );
  DFFPOSX1 ram_reg_160__1_ ( .D(n6998), .CLK(clk), .Q(ram[2561]) );
  DFFPOSX1 ram_reg_160__0_ ( .D(n6997), .CLK(clk), .Q(ram[2560]) );
  DFFPOSX1 ram_reg_159__15_ ( .D(n6996), .CLK(clk), .Q(ram[2559]) );
  DFFPOSX1 ram_reg_159__14_ ( .D(n6995), .CLK(clk), .Q(ram[2558]) );
  DFFPOSX1 ram_reg_159__13_ ( .D(n6994), .CLK(clk), .Q(ram[2557]) );
  DFFPOSX1 ram_reg_159__12_ ( .D(n6993), .CLK(clk), .Q(ram[2556]) );
  DFFPOSX1 ram_reg_159__11_ ( .D(n6992), .CLK(clk), .Q(ram[2555]) );
  DFFPOSX1 ram_reg_159__10_ ( .D(n6991), .CLK(clk), .Q(ram[2554]) );
  DFFPOSX1 ram_reg_159__9_ ( .D(n6990), .CLK(clk), .Q(ram[2553]) );
  DFFPOSX1 ram_reg_159__8_ ( .D(n6989), .CLK(clk), .Q(ram[2552]) );
  DFFPOSX1 ram_reg_159__7_ ( .D(n6988), .CLK(clk), .Q(ram[2551]) );
  DFFPOSX1 ram_reg_159__6_ ( .D(n6987), .CLK(clk), .Q(ram[2550]) );
  DFFPOSX1 ram_reg_159__5_ ( .D(n6986), .CLK(clk), .Q(ram[2549]) );
  DFFPOSX1 ram_reg_159__4_ ( .D(n6985), .CLK(clk), .Q(ram[2548]) );
  DFFPOSX1 ram_reg_159__3_ ( .D(n6984), .CLK(clk), .Q(ram[2547]) );
  DFFPOSX1 ram_reg_159__2_ ( .D(n6983), .CLK(clk), .Q(ram[2546]) );
  DFFPOSX1 ram_reg_159__1_ ( .D(n6982), .CLK(clk), .Q(ram[2545]) );
  DFFPOSX1 ram_reg_159__0_ ( .D(n6981), .CLK(clk), .Q(ram[2544]) );
  DFFPOSX1 ram_reg_158__15_ ( .D(n6980), .CLK(clk), .Q(ram[2543]) );
  DFFPOSX1 ram_reg_158__14_ ( .D(n6979), .CLK(clk), .Q(ram[2542]) );
  DFFPOSX1 ram_reg_158__13_ ( .D(n6978), .CLK(clk), .Q(ram[2541]) );
  DFFPOSX1 ram_reg_158__12_ ( .D(n6977), .CLK(clk), .Q(ram[2540]) );
  DFFPOSX1 ram_reg_158__11_ ( .D(n6976), .CLK(clk), .Q(ram[2539]) );
  DFFPOSX1 ram_reg_158__10_ ( .D(n6975), .CLK(clk), .Q(ram[2538]) );
  DFFPOSX1 ram_reg_158__9_ ( .D(n6974), .CLK(clk), .Q(ram[2537]) );
  DFFPOSX1 ram_reg_158__8_ ( .D(n6973), .CLK(clk), .Q(ram[2536]) );
  DFFPOSX1 ram_reg_158__7_ ( .D(n6972), .CLK(clk), .Q(ram[2535]) );
  DFFPOSX1 ram_reg_158__6_ ( .D(n6971), .CLK(clk), .Q(ram[2534]) );
  DFFPOSX1 ram_reg_158__5_ ( .D(n6970), .CLK(clk), .Q(ram[2533]) );
  DFFPOSX1 ram_reg_158__4_ ( .D(n6969), .CLK(clk), .Q(ram[2532]) );
  DFFPOSX1 ram_reg_158__3_ ( .D(n6968), .CLK(clk), .Q(ram[2531]) );
  DFFPOSX1 ram_reg_158__2_ ( .D(n6967), .CLK(clk), .Q(ram[2530]) );
  DFFPOSX1 ram_reg_158__1_ ( .D(n6966), .CLK(clk), .Q(ram[2529]) );
  DFFPOSX1 ram_reg_158__0_ ( .D(n6965), .CLK(clk), .Q(ram[2528]) );
  DFFPOSX1 ram_reg_157__15_ ( .D(n6964), .CLK(clk), .Q(ram[2527]) );
  DFFPOSX1 ram_reg_157__14_ ( .D(n6963), .CLK(clk), .Q(ram[2526]) );
  DFFPOSX1 ram_reg_157__13_ ( .D(n6962), .CLK(clk), .Q(ram[2525]) );
  DFFPOSX1 ram_reg_157__12_ ( .D(n6961), .CLK(clk), .Q(ram[2524]) );
  DFFPOSX1 ram_reg_157__11_ ( .D(n6960), .CLK(clk), .Q(ram[2523]) );
  DFFPOSX1 ram_reg_157__10_ ( .D(n6959), .CLK(clk), .Q(ram[2522]) );
  DFFPOSX1 ram_reg_157__9_ ( .D(n6958), .CLK(clk), .Q(ram[2521]) );
  DFFPOSX1 ram_reg_157__8_ ( .D(n6957), .CLK(clk), .Q(ram[2520]) );
  DFFPOSX1 ram_reg_157__7_ ( .D(n6956), .CLK(clk), .Q(ram[2519]) );
  DFFPOSX1 ram_reg_157__6_ ( .D(n6955), .CLK(clk), .Q(ram[2518]) );
  DFFPOSX1 ram_reg_157__5_ ( .D(n6954), .CLK(clk), .Q(ram[2517]) );
  DFFPOSX1 ram_reg_157__4_ ( .D(n6953), .CLK(clk), .Q(ram[2516]) );
  DFFPOSX1 ram_reg_157__3_ ( .D(n6952), .CLK(clk), .Q(ram[2515]) );
  DFFPOSX1 ram_reg_157__2_ ( .D(n6951), .CLK(clk), .Q(ram[2514]) );
  DFFPOSX1 ram_reg_157__1_ ( .D(n6950), .CLK(clk), .Q(ram[2513]) );
  DFFPOSX1 ram_reg_157__0_ ( .D(n6949), .CLK(clk), .Q(ram[2512]) );
  DFFPOSX1 ram_reg_156__15_ ( .D(n6948), .CLK(clk), .Q(ram[2511]) );
  DFFPOSX1 ram_reg_156__14_ ( .D(n6947), .CLK(clk), .Q(ram[2510]) );
  DFFPOSX1 ram_reg_156__13_ ( .D(n6946), .CLK(clk), .Q(ram[2509]) );
  DFFPOSX1 ram_reg_156__12_ ( .D(n6945), .CLK(clk), .Q(ram[2508]) );
  DFFPOSX1 ram_reg_156__11_ ( .D(n6944), .CLK(clk), .Q(ram[2507]) );
  DFFPOSX1 ram_reg_156__10_ ( .D(n6943), .CLK(clk), .Q(ram[2506]) );
  DFFPOSX1 ram_reg_156__9_ ( .D(n6942), .CLK(clk), .Q(ram[2505]) );
  DFFPOSX1 ram_reg_156__8_ ( .D(n6941), .CLK(clk), .Q(ram[2504]) );
  DFFPOSX1 ram_reg_156__7_ ( .D(n6940), .CLK(clk), .Q(ram[2503]) );
  DFFPOSX1 ram_reg_156__6_ ( .D(n6939), .CLK(clk), .Q(ram[2502]) );
  DFFPOSX1 ram_reg_156__5_ ( .D(n6938), .CLK(clk), .Q(ram[2501]) );
  DFFPOSX1 ram_reg_156__4_ ( .D(n6937), .CLK(clk), .Q(ram[2500]) );
  DFFPOSX1 ram_reg_156__3_ ( .D(n6936), .CLK(clk), .Q(ram[2499]) );
  DFFPOSX1 ram_reg_156__2_ ( .D(n6935), .CLK(clk), .Q(ram[2498]) );
  DFFPOSX1 ram_reg_156__1_ ( .D(n6934), .CLK(clk), .Q(ram[2497]) );
  DFFPOSX1 ram_reg_156__0_ ( .D(n6933), .CLK(clk), .Q(ram[2496]) );
  DFFPOSX1 ram_reg_155__15_ ( .D(n6932), .CLK(clk), .Q(ram[2495]) );
  DFFPOSX1 ram_reg_155__14_ ( .D(n6931), .CLK(clk), .Q(ram[2494]) );
  DFFPOSX1 ram_reg_155__13_ ( .D(n6930), .CLK(clk), .Q(ram[2493]) );
  DFFPOSX1 ram_reg_155__12_ ( .D(n6929), .CLK(clk), .Q(ram[2492]) );
  DFFPOSX1 ram_reg_155__11_ ( .D(n6928), .CLK(clk), .Q(ram[2491]) );
  DFFPOSX1 ram_reg_155__10_ ( .D(n6927), .CLK(clk), .Q(ram[2490]) );
  DFFPOSX1 ram_reg_155__9_ ( .D(n6926), .CLK(clk), .Q(ram[2489]) );
  DFFPOSX1 ram_reg_155__8_ ( .D(n6925), .CLK(clk), .Q(ram[2488]) );
  DFFPOSX1 ram_reg_155__7_ ( .D(n6924), .CLK(clk), .Q(ram[2487]) );
  DFFPOSX1 ram_reg_155__6_ ( .D(n6923), .CLK(clk), .Q(ram[2486]) );
  DFFPOSX1 ram_reg_155__5_ ( .D(n6922), .CLK(clk), .Q(ram[2485]) );
  DFFPOSX1 ram_reg_155__4_ ( .D(n6921), .CLK(clk), .Q(ram[2484]) );
  DFFPOSX1 ram_reg_155__3_ ( .D(n6920), .CLK(clk), .Q(ram[2483]) );
  DFFPOSX1 ram_reg_155__2_ ( .D(n6919), .CLK(clk), .Q(ram[2482]) );
  DFFPOSX1 ram_reg_155__1_ ( .D(n6918), .CLK(clk), .Q(ram[2481]) );
  DFFPOSX1 ram_reg_155__0_ ( .D(n6917), .CLK(clk), .Q(ram[2480]) );
  DFFPOSX1 ram_reg_154__15_ ( .D(n6916), .CLK(clk), .Q(ram[2479]) );
  DFFPOSX1 ram_reg_154__14_ ( .D(n6915), .CLK(clk), .Q(ram[2478]) );
  DFFPOSX1 ram_reg_154__13_ ( .D(n6914), .CLK(clk), .Q(ram[2477]) );
  DFFPOSX1 ram_reg_154__12_ ( .D(n6913), .CLK(clk), .Q(ram[2476]) );
  DFFPOSX1 ram_reg_154__11_ ( .D(n6912), .CLK(clk), .Q(ram[2475]) );
  DFFPOSX1 ram_reg_154__10_ ( .D(n6911), .CLK(clk), .Q(ram[2474]) );
  DFFPOSX1 ram_reg_154__9_ ( .D(n6910), .CLK(clk), .Q(ram[2473]) );
  DFFPOSX1 ram_reg_154__8_ ( .D(n6909), .CLK(clk), .Q(ram[2472]) );
  DFFPOSX1 ram_reg_154__7_ ( .D(n6908), .CLK(clk), .Q(ram[2471]) );
  DFFPOSX1 ram_reg_154__6_ ( .D(n6907), .CLK(clk), .Q(ram[2470]) );
  DFFPOSX1 ram_reg_154__5_ ( .D(n6906), .CLK(clk), .Q(ram[2469]) );
  DFFPOSX1 ram_reg_154__4_ ( .D(n6905), .CLK(clk), .Q(ram[2468]) );
  DFFPOSX1 ram_reg_154__3_ ( .D(n6904), .CLK(clk), .Q(ram[2467]) );
  DFFPOSX1 ram_reg_154__2_ ( .D(n6903), .CLK(clk), .Q(ram[2466]) );
  DFFPOSX1 ram_reg_154__1_ ( .D(n6902), .CLK(clk), .Q(ram[2465]) );
  DFFPOSX1 ram_reg_154__0_ ( .D(n6901), .CLK(clk), .Q(ram[2464]) );
  DFFPOSX1 ram_reg_153__15_ ( .D(n6900), .CLK(clk), .Q(ram[2463]) );
  DFFPOSX1 ram_reg_153__14_ ( .D(n6899), .CLK(clk), .Q(ram[2462]) );
  DFFPOSX1 ram_reg_153__13_ ( .D(n6898), .CLK(clk), .Q(ram[2461]) );
  DFFPOSX1 ram_reg_153__12_ ( .D(n6897), .CLK(clk), .Q(ram[2460]) );
  DFFPOSX1 ram_reg_153__11_ ( .D(n6896), .CLK(clk), .Q(ram[2459]) );
  DFFPOSX1 ram_reg_153__10_ ( .D(n6895), .CLK(clk), .Q(ram[2458]) );
  DFFPOSX1 ram_reg_153__9_ ( .D(n6894), .CLK(clk), .Q(ram[2457]) );
  DFFPOSX1 ram_reg_153__8_ ( .D(n6893), .CLK(clk), .Q(ram[2456]) );
  DFFPOSX1 ram_reg_153__7_ ( .D(n6892), .CLK(clk), .Q(ram[2455]) );
  DFFPOSX1 ram_reg_153__6_ ( .D(n6891), .CLK(clk), .Q(ram[2454]) );
  DFFPOSX1 ram_reg_153__5_ ( .D(n6890), .CLK(clk), .Q(ram[2453]) );
  DFFPOSX1 ram_reg_153__4_ ( .D(n6889), .CLK(clk), .Q(ram[2452]) );
  DFFPOSX1 ram_reg_153__3_ ( .D(n6888), .CLK(clk), .Q(ram[2451]) );
  DFFPOSX1 ram_reg_153__2_ ( .D(n6887), .CLK(clk), .Q(ram[2450]) );
  DFFPOSX1 ram_reg_153__1_ ( .D(n6886), .CLK(clk), .Q(ram[2449]) );
  DFFPOSX1 ram_reg_153__0_ ( .D(n6885), .CLK(clk), .Q(ram[2448]) );
  DFFPOSX1 ram_reg_152__15_ ( .D(n6884), .CLK(clk), .Q(ram[2447]) );
  DFFPOSX1 ram_reg_152__14_ ( .D(n6883), .CLK(clk), .Q(ram[2446]) );
  DFFPOSX1 ram_reg_152__13_ ( .D(n6882), .CLK(clk), .Q(ram[2445]) );
  DFFPOSX1 ram_reg_152__12_ ( .D(n6881), .CLK(clk), .Q(ram[2444]) );
  DFFPOSX1 ram_reg_152__11_ ( .D(n6880), .CLK(clk), .Q(ram[2443]) );
  DFFPOSX1 ram_reg_152__10_ ( .D(n6879), .CLK(clk), .Q(ram[2442]) );
  DFFPOSX1 ram_reg_152__9_ ( .D(n6878), .CLK(clk), .Q(ram[2441]) );
  DFFPOSX1 ram_reg_152__8_ ( .D(n6877), .CLK(clk), .Q(ram[2440]) );
  DFFPOSX1 ram_reg_152__7_ ( .D(n6876), .CLK(clk), .Q(ram[2439]) );
  DFFPOSX1 ram_reg_152__6_ ( .D(n6875), .CLK(clk), .Q(ram[2438]) );
  DFFPOSX1 ram_reg_152__5_ ( .D(n6874), .CLK(clk), .Q(ram[2437]) );
  DFFPOSX1 ram_reg_152__4_ ( .D(n6873), .CLK(clk), .Q(ram[2436]) );
  DFFPOSX1 ram_reg_152__3_ ( .D(n6872), .CLK(clk), .Q(ram[2435]) );
  DFFPOSX1 ram_reg_152__2_ ( .D(n6871), .CLK(clk), .Q(ram[2434]) );
  DFFPOSX1 ram_reg_152__1_ ( .D(n6870), .CLK(clk), .Q(ram[2433]) );
  DFFPOSX1 ram_reg_152__0_ ( .D(n6869), .CLK(clk), .Q(ram[2432]) );
  DFFPOSX1 ram_reg_151__15_ ( .D(n6868), .CLK(clk), .Q(ram[2431]) );
  DFFPOSX1 ram_reg_151__14_ ( .D(n6867), .CLK(clk), .Q(ram[2430]) );
  DFFPOSX1 ram_reg_151__13_ ( .D(n6866), .CLK(clk), .Q(ram[2429]) );
  DFFPOSX1 ram_reg_151__12_ ( .D(n6865), .CLK(clk), .Q(ram[2428]) );
  DFFPOSX1 ram_reg_151__11_ ( .D(n6864), .CLK(clk), .Q(ram[2427]) );
  DFFPOSX1 ram_reg_151__10_ ( .D(n6863), .CLK(clk), .Q(ram[2426]) );
  DFFPOSX1 ram_reg_151__9_ ( .D(n6862), .CLK(clk), .Q(ram[2425]) );
  DFFPOSX1 ram_reg_151__8_ ( .D(n6861), .CLK(clk), .Q(ram[2424]) );
  DFFPOSX1 ram_reg_151__7_ ( .D(n6860), .CLK(clk), .Q(ram[2423]) );
  DFFPOSX1 ram_reg_151__6_ ( .D(n6859), .CLK(clk), .Q(ram[2422]) );
  DFFPOSX1 ram_reg_151__5_ ( .D(n6858), .CLK(clk), .Q(ram[2421]) );
  DFFPOSX1 ram_reg_151__4_ ( .D(n6857), .CLK(clk), .Q(ram[2420]) );
  DFFPOSX1 ram_reg_151__3_ ( .D(n6856), .CLK(clk), .Q(ram[2419]) );
  DFFPOSX1 ram_reg_151__2_ ( .D(n6855), .CLK(clk), .Q(ram[2418]) );
  DFFPOSX1 ram_reg_151__1_ ( .D(n6854), .CLK(clk), .Q(ram[2417]) );
  DFFPOSX1 ram_reg_151__0_ ( .D(n6853), .CLK(clk), .Q(ram[2416]) );
  DFFPOSX1 ram_reg_150__15_ ( .D(n6852), .CLK(clk), .Q(ram[2415]) );
  DFFPOSX1 ram_reg_150__14_ ( .D(n6851), .CLK(clk), .Q(ram[2414]) );
  DFFPOSX1 ram_reg_150__13_ ( .D(n6850), .CLK(clk), .Q(ram[2413]) );
  DFFPOSX1 ram_reg_150__12_ ( .D(n6849), .CLK(clk), .Q(ram[2412]) );
  DFFPOSX1 ram_reg_150__11_ ( .D(n6848), .CLK(clk), .Q(ram[2411]) );
  DFFPOSX1 ram_reg_150__10_ ( .D(n6847), .CLK(clk), .Q(ram[2410]) );
  DFFPOSX1 ram_reg_150__9_ ( .D(n6846), .CLK(clk), .Q(ram[2409]) );
  DFFPOSX1 ram_reg_150__8_ ( .D(n6845), .CLK(clk), .Q(ram[2408]) );
  DFFPOSX1 ram_reg_150__7_ ( .D(n6844), .CLK(clk), .Q(ram[2407]) );
  DFFPOSX1 ram_reg_150__6_ ( .D(n6843), .CLK(clk), .Q(ram[2406]) );
  DFFPOSX1 ram_reg_150__5_ ( .D(n6842), .CLK(clk), .Q(ram[2405]) );
  DFFPOSX1 ram_reg_150__4_ ( .D(n6841), .CLK(clk), .Q(ram[2404]) );
  DFFPOSX1 ram_reg_150__3_ ( .D(n6840), .CLK(clk), .Q(ram[2403]) );
  DFFPOSX1 ram_reg_150__2_ ( .D(n6839), .CLK(clk), .Q(ram[2402]) );
  DFFPOSX1 ram_reg_150__1_ ( .D(n6838), .CLK(clk), .Q(ram[2401]) );
  DFFPOSX1 ram_reg_150__0_ ( .D(n6837), .CLK(clk), .Q(ram[2400]) );
  DFFPOSX1 ram_reg_149__15_ ( .D(n6836), .CLK(clk), .Q(ram[2399]) );
  DFFPOSX1 ram_reg_149__14_ ( .D(n6835), .CLK(clk), .Q(ram[2398]) );
  DFFPOSX1 ram_reg_149__13_ ( .D(n6834), .CLK(clk), .Q(ram[2397]) );
  DFFPOSX1 ram_reg_149__12_ ( .D(n6833), .CLK(clk), .Q(ram[2396]) );
  DFFPOSX1 ram_reg_149__11_ ( .D(n6832), .CLK(clk), .Q(ram[2395]) );
  DFFPOSX1 ram_reg_149__10_ ( .D(n6831), .CLK(clk), .Q(ram[2394]) );
  DFFPOSX1 ram_reg_149__9_ ( .D(n6830), .CLK(clk), .Q(ram[2393]) );
  DFFPOSX1 ram_reg_149__8_ ( .D(n6829), .CLK(clk), .Q(ram[2392]) );
  DFFPOSX1 ram_reg_149__7_ ( .D(n6828), .CLK(clk), .Q(ram[2391]) );
  DFFPOSX1 ram_reg_149__6_ ( .D(n6827), .CLK(clk), .Q(ram[2390]) );
  DFFPOSX1 ram_reg_149__5_ ( .D(n6826), .CLK(clk), .Q(ram[2389]) );
  DFFPOSX1 ram_reg_149__4_ ( .D(n6825), .CLK(clk), .Q(ram[2388]) );
  DFFPOSX1 ram_reg_149__3_ ( .D(n6824), .CLK(clk), .Q(ram[2387]) );
  DFFPOSX1 ram_reg_149__2_ ( .D(n6823), .CLK(clk), .Q(ram[2386]) );
  DFFPOSX1 ram_reg_149__1_ ( .D(n6822), .CLK(clk), .Q(ram[2385]) );
  DFFPOSX1 ram_reg_149__0_ ( .D(n6821), .CLK(clk), .Q(ram[2384]) );
  DFFPOSX1 ram_reg_148__15_ ( .D(n6820), .CLK(clk), .Q(ram[2383]) );
  DFFPOSX1 ram_reg_148__14_ ( .D(n6819), .CLK(clk), .Q(ram[2382]) );
  DFFPOSX1 ram_reg_148__13_ ( .D(n6818), .CLK(clk), .Q(ram[2381]) );
  DFFPOSX1 ram_reg_148__12_ ( .D(n6817), .CLK(clk), .Q(ram[2380]) );
  DFFPOSX1 ram_reg_148__11_ ( .D(n6816), .CLK(clk), .Q(ram[2379]) );
  DFFPOSX1 ram_reg_148__10_ ( .D(n6815), .CLK(clk), .Q(ram[2378]) );
  DFFPOSX1 ram_reg_148__9_ ( .D(n6814), .CLK(clk), .Q(ram[2377]) );
  DFFPOSX1 ram_reg_148__8_ ( .D(n6813), .CLK(clk), .Q(ram[2376]) );
  DFFPOSX1 ram_reg_148__7_ ( .D(n6812), .CLK(clk), .Q(ram[2375]) );
  DFFPOSX1 ram_reg_148__6_ ( .D(n6811), .CLK(clk), .Q(ram[2374]) );
  DFFPOSX1 ram_reg_148__5_ ( .D(n6810), .CLK(clk), .Q(ram[2373]) );
  DFFPOSX1 ram_reg_148__4_ ( .D(n6809), .CLK(clk), .Q(ram[2372]) );
  DFFPOSX1 ram_reg_148__3_ ( .D(n6808), .CLK(clk), .Q(ram[2371]) );
  DFFPOSX1 ram_reg_148__2_ ( .D(n6807), .CLK(clk), .Q(ram[2370]) );
  DFFPOSX1 ram_reg_148__1_ ( .D(n6806), .CLK(clk), .Q(ram[2369]) );
  DFFPOSX1 ram_reg_148__0_ ( .D(n6805), .CLK(clk), .Q(ram[2368]) );
  DFFPOSX1 ram_reg_147__15_ ( .D(n6804), .CLK(clk), .Q(ram[2367]) );
  DFFPOSX1 ram_reg_147__14_ ( .D(n6803), .CLK(clk), .Q(ram[2366]) );
  DFFPOSX1 ram_reg_147__13_ ( .D(n6802), .CLK(clk), .Q(ram[2365]) );
  DFFPOSX1 ram_reg_147__12_ ( .D(n6801), .CLK(clk), .Q(ram[2364]) );
  DFFPOSX1 ram_reg_147__11_ ( .D(n6800), .CLK(clk), .Q(ram[2363]) );
  DFFPOSX1 ram_reg_147__10_ ( .D(n6799), .CLK(clk), .Q(ram[2362]) );
  DFFPOSX1 ram_reg_147__9_ ( .D(n6798), .CLK(clk), .Q(ram[2361]) );
  DFFPOSX1 ram_reg_147__8_ ( .D(n6797), .CLK(clk), .Q(ram[2360]) );
  DFFPOSX1 ram_reg_147__7_ ( .D(n6796), .CLK(clk), .Q(ram[2359]) );
  DFFPOSX1 ram_reg_147__6_ ( .D(n6795), .CLK(clk), .Q(ram[2358]) );
  DFFPOSX1 ram_reg_147__5_ ( .D(n6794), .CLK(clk), .Q(ram[2357]) );
  DFFPOSX1 ram_reg_147__4_ ( .D(n6793), .CLK(clk), .Q(ram[2356]) );
  DFFPOSX1 ram_reg_147__3_ ( .D(n6792), .CLK(clk), .Q(ram[2355]) );
  DFFPOSX1 ram_reg_147__2_ ( .D(n6791), .CLK(clk), .Q(ram[2354]) );
  DFFPOSX1 ram_reg_147__1_ ( .D(n6790), .CLK(clk), .Q(ram[2353]) );
  DFFPOSX1 ram_reg_147__0_ ( .D(n6789), .CLK(clk), .Q(ram[2352]) );
  DFFPOSX1 ram_reg_146__15_ ( .D(n6788), .CLK(clk), .Q(ram[2351]) );
  DFFPOSX1 ram_reg_146__14_ ( .D(n6787), .CLK(clk), .Q(ram[2350]) );
  DFFPOSX1 ram_reg_146__13_ ( .D(n6786), .CLK(clk), .Q(ram[2349]) );
  DFFPOSX1 ram_reg_146__12_ ( .D(n6785), .CLK(clk), .Q(ram[2348]) );
  DFFPOSX1 ram_reg_146__11_ ( .D(n6784), .CLK(clk), .Q(ram[2347]) );
  DFFPOSX1 ram_reg_146__10_ ( .D(n6783), .CLK(clk), .Q(ram[2346]) );
  DFFPOSX1 ram_reg_146__9_ ( .D(n6782), .CLK(clk), .Q(ram[2345]) );
  DFFPOSX1 ram_reg_146__8_ ( .D(n6781), .CLK(clk), .Q(ram[2344]) );
  DFFPOSX1 ram_reg_146__7_ ( .D(n6780), .CLK(clk), .Q(ram[2343]) );
  DFFPOSX1 ram_reg_146__6_ ( .D(n6779), .CLK(clk), .Q(ram[2342]) );
  DFFPOSX1 ram_reg_146__5_ ( .D(n6778), .CLK(clk), .Q(ram[2341]) );
  DFFPOSX1 ram_reg_146__4_ ( .D(n6777), .CLK(clk), .Q(ram[2340]) );
  DFFPOSX1 ram_reg_146__3_ ( .D(n6776), .CLK(clk), .Q(ram[2339]) );
  DFFPOSX1 ram_reg_146__2_ ( .D(n6775), .CLK(clk), .Q(ram[2338]) );
  DFFPOSX1 ram_reg_146__1_ ( .D(n6774), .CLK(clk), .Q(ram[2337]) );
  DFFPOSX1 ram_reg_146__0_ ( .D(n6773), .CLK(clk), .Q(ram[2336]) );
  DFFPOSX1 ram_reg_145__15_ ( .D(n6772), .CLK(clk), .Q(ram[2335]) );
  DFFPOSX1 ram_reg_145__14_ ( .D(n6771), .CLK(clk), .Q(ram[2334]) );
  DFFPOSX1 ram_reg_145__13_ ( .D(n6770), .CLK(clk), .Q(ram[2333]) );
  DFFPOSX1 ram_reg_145__12_ ( .D(n6769), .CLK(clk), .Q(ram[2332]) );
  DFFPOSX1 ram_reg_145__11_ ( .D(n6768), .CLK(clk), .Q(ram[2331]) );
  DFFPOSX1 ram_reg_145__10_ ( .D(n6767), .CLK(clk), .Q(ram[2330]) );
  DFFPOSX1 ram_reg_145__9_ ( .D(n6766), .CLK(clk), .Q(ram[2329]) );
  DFFPOSX1 ram_reg_145__8_ ( .D(n6765), .CLK(clk), .Q(ram[2328]) );
  DFFPOSX1 ram_reg_145__7_ ( .D(n6764), .CLK(clk), .Q(ram[2327]) );
  DFFPOSX1 ram_reg_145__6_ ( .D(n6763), .CLK(clk), .Q(ram[2326]) );
  DFFPOSX1 ram_reg_145__5_ ( .D(n6762), .CLK(clk), .Q(ram[2325]) );
  DFFPOSX1 ram_reg_145__4_ ( .D(n6761), .CLK(clk), .Q(ram[2324]) );
  DFFPOSX1 ram_reg_145__3_ ( .D(n6760), .CLK(clk), .Q(ram[2323]) );
  DFFPOSX1 ram_reg_145__2_ ( .D(n6759), .CLK(clk), .Q(ram[2322]) );
  DFFPOSX1 ram_reg_145__1_ ( .D(n6758), .CLK(clk), .Q(ram[2321]) );
  DFFPOSX1 ram_reg_145__0_ ( .D(n6757), .CLK(clk), .Q(ram[2320]) );
  DFFPOSX1 ram_reg_144__15_ ( .D(n6756), .CLK(clk), .Q(ram[2319]) );
  DFFPOSX1 ram_reg_144__14_ ( .D(n6755), .CLK(clk), .Q(ram[2318]) );
  DFFPOSX1 ram_reg_144__13_ ( .D(n6754), .CLK(clk), .Q(ram[2317]) );
  DFFPOSX1 ram_reg_144__12_ ( .D(n6753), .CLK(clk), .Q(ram[2316]) );
  DFFPOSX1 ram_reg_144__11_ ( .D(n6752), .CLK(clk), .Q(ram[2315]) );
  DFFPOSX1 ram_reg_144__10_ ( .D(n6751), .CLK(clk), .Q(ram[2314]) );
  DFFPOSX1 ram_reg_144__9_ ( .D(n6750), .CLK(clk), .Q(ram[2313]) );
  DFFPOSX1 ram_reg_144__8_ ( .D(n6749), .CLK(clk), .Q(ram[2312]) );
  DFFPOSX1 ram_reg_144__7_ ( .D(n6748), .CLK(clk), .Q(ram[2311]) );
  DFFPOSX1 ram_reg_144__6_ ( .D(n6747), .CLK(clk), .Q(ram[2310]) );
  DFFPOSX1 ram_reg_144__5_ ( .D(n6746), .CLK(clk), .Q(ram[2309]) );
  DFFPOSX1 ram_reg_144__4_ ( .D(n6745), .CLK(clk), .Q(ram[2308]) );
  DFFPOSX1 ram_reg_144__3_ ( .D(n6744), .CLK(clk), .Q(ram[2307]) );
  DFFPOSX1 ram_reg_144__2_ ( .D(n6743), .CLK(clk), .Q(ram[2306]) );
  DFFPOSX1 ram_reg_144__1_ ( .D(n6742), .CLK(clk), .Q(ram[2305]) );
  DFFPOSX1 ram_reg_144__0_ ( .D(n6741), .CLK(clk), .Q(ram[2304]) );
  DFFPOSX1 ram_reg_143__15_ ( .D(n6740), .CLK(clk), .Q(ram[2303]) );
  DFFPOSX1 ram_reg_143__14_ ( .D(n6739), .CLK(clk), .Q(ram[2302]) );
  DFFPOSX1 ram_reg_143__13_ ( .D(n6738), .CLK(clk), .Q(ram[2301]) );
  DFFPOSX1 ram_reg_143__12_ ( .D(n6737), .CLK(clk), .Q(ram[2300]) );
  DFFPOSX1 ram_reg_143__11_ ( .D(n6736), .CLK(clk), .Q(ram[2299]) );
  DFFPOSX1 ram_reg_143__10_ ( .D(n6735), .CLK(clk), .Q(ram[2298]) );
  DFFPOSX1 ram_reg_143__9_ ( .D(n6734), .CLK(clk), .Q(ram[2297]) );
  DFFPOSX1 ram_reg_143__8_ ( .D(n6733), .CLK(clk), .Q(ram[2296]) );
  DFFPOSX1 ram_reg_143__7_ ( .D(n6732), .CLK(clk), .Q(ram[2295]) );
  DFFPOSX1 ram_reg_143__6_ ( .D(n6731), .CLK(clk), .Q(ram[2294]) );
  DFFPOSX1 ram_reg_143__5_ ( .D(n6730), .CLK(clk), .Q(ram[2293]) );
  DFFPOSX1 ram_reg_143__4_ ( .D(n6729), .CLK(clk), .Q(ram[2292]) );
  DFFPOSX1 ram_reg_143__3_ ( .D(n6728), .CLK(clk), .Q(ram[2291]) );
  DFFPOSX1 ram_reg_143__2_ ( .D(n6727), .CLK(clk), .Q(ram[2290]) );
  DFFPOSX1 ram_reg_143__1_ ( .D(n6726), .CLK(clk), .Q(ram[2289]) );
  DFFPOSX1 ram_reg_143__0_ ( .D(n6725), .CLK(clk), .Q(ram[2288]) );
  DFFPOSX1 ram_reg_142__15_ ( .D(n6724), .CLK(clk), .Q(ram[2287]) );
  DFFPOSX1 ram_reg_142__14_ ( .D(n6723), .CLK(clk), .Q(ram[2286]) );
  DFFPOSX1 ram_reg_142__13_ ( .D(n6722), .CLK(clk), .Q(ram[2285]) );
  DFFPOSX1 ram_reg_142__12_ ( .D(n6721), .CLK(clk), .Q(ram[2284]) );
  DFFPOSX1 ram_reg_142__11_ ( .D(n6720), .CLK(clk), .Q(ram[2283]) );
  DFFPOSX1 ram_reg_142__10_ ( .D(n6719), .CLK(clk), .Q(ram[2282]) );
  DFFPOSX1 ram_reg_142__9_ ( .D(n6718), .CLK(clk), .Q(ram[2281]) );
  DFFPOSX1 ram_reg_142__8_ ( .D(n6717), .CLK(clk), .Q(ram[2280]) );
  DFFPOSX1 ram_reg_142__7_ ( .D(n6716), .CLK(clk), .Q(ram[2279]) );
  DFFPOSX1 ram_reg_142__6_ ( .D(n6715), .CLK(clk), .Q(ram[2278]) );
  DFFPOSX1 ram_reg_142__5_ ( .D(n6714), .CLK(clk), .Q(ram[2277]) );
  DFFPOSX1 ram_reg_142__4_ ( .D(n6713), .CLK(clk), .Q(ram[2276]) );
  DFFPOSX1 ram_reg_142__3_ ( .D(n6712), .CLK(clk), .Q(ram[2275]) );
  DFFPOSX1 ram_reg_142__2_ ( .D(n6711), .CLK(clk), .Q(ram[2274]) );
  DFFPOSX1 ram_reg_142__1_ ( .D(n6710), .CLK(clk), .Q(ram[2273]) );
  DFFPOSX1 ram_reg_142__0_ ( .D(n6709), .CLK(clk), .Q(ram[2272]) );
  DFFPOSX1 ram_reg_141__15_ ( .D(n6708), .CLK(clk), .Q(ram[2271]) );
  DFFPOSX1 ram_reg_141__14_ ( .D(n6707), .CLK(clk), .Q(ram[2270]) );
  DFFPOSX1 ram_reg_141__13_ ( .D(n6706), .CLK(clk), .Q(ram[2269]) );
  DFFPOSX1 ram_reg_141__12_ ( .D(n6705), .CLK(clk), .Q(ram[2268]) );
  DFFPOSX1 ram_reg_141__11_ ( .D(n6704), .CLK(clk), .Q(ram[2267]) );
  DFFPOSX1 ram_reg_141__10_ ( .D(n6703), .CLK(clk), .Q(ram[2266]) );
  DFFPOSX1 ram_reg_141__9_ ( .D(n6702), .CLK(clk), .Q(ram[2265]) );
  DFFPOSX1 ram_reg_141__8_ ( .D(n6701), .CLK(clk), .Q(ram[2264]) );
  DFFPOSX1 ram_reg_141__7_ ( .D(n6700), .CLK(clk), .Q(ram[2263]) );
  DFFPOSX1 ram_reg_141__6_ ( .D(n6699), .CLK(clk), .Q(ram[2262]) );
  DFFPOSX1 ram_reg_141__5_ ( .D(n6698), .CLK(clk), .Q(ram[2261]) );
  DFFPOSX1 ram_reg_141__4_ ( .D(n6697), .CLK(clk), .Q(ram[2260]) );
  DFFPOSX1 ram_reg_141__3_ ( .D(n6696), .CLK(clk), .Q(ram[2259]) );
  DFFPOSX1 ram_reg_141__2_ ( .D(n6695), .CLK(clk), .Q(ram[2258]) );
  DFFPOSX1 ram_reg_141__1_ ( .D(n6694), .CLK(clk), .Q(ram[2257]) );
  DFFPOSX1 ram_reg_141__0_ ( .D(n6693), .CLK(clk), .Q(ram[2256]) );
  DFFPOSX1 ram_reg_140__15_ ( .D(n6692), .CLK(clk), .Q(ram[2255]) );
  DFFPOSX1 ram_reg_140__14_ ( .D(n6691), .CLK(clk), .Q(ram[2254]) );
  DFFPOSX1 ram_reg_140__13_ ( .D(n6690), .CLK(clk), .Q(ram[2253]) );
  DFFPOSX1 ram_reg_140__12_ ( .D(n6689), .CLK(clk), .Q(ram[2252]) );
  DFFPOSX1 ram_reg_140__11_ ( .D(n6688), .CLK(clk), .Q(ram[2251]) );
  DFFPOSX1 ram_reg_140__10_ ( .D(n6687), .CLK(clk), .Q(ram[2250]) );
  DFFPOSX1 ram_reg_140__9_ ( .D(n6686), .CLK(clk), .Q(ram[2249]) );
  DFFPOSX1 ram_reg_140__8_ ( .D(n6685), .CLK(clk), .Q(ram[2248]) );
  DFFPOSX1 ram_reg_140__7_ ( .D(n6684), .CLK(clk), .Q(ram[2247]) );
  DFFPOSX1 ram_reg_140__6_ ( .D(n6683), .CLK(clk), .Q(ram[2246]) );
  DFFPOSX1 ram_reg_140__5_ ( .D(n6682), .CLK(clk), .Q(ram[2245]) );
  DFFPOSX1 ram_reg_140__4_ ( .D(n6681), .CLK(clk), .Q(ram[2244]) );
  DFFPOSX1 ram_reg_140__3_ ( .D(n6680), .CLK(clk), .Q(ram[2243]) );
  DFFPOSX1 ram_reg_140__2_ ( .D(n6679), .CLK(clk), .Q(ram[2242]) );
  DFFPOSX1 ram_reg_140__1_ ( .D(n6678), .CLK(clk), .Q(ram[2241]) );
  DFFPOSX1 ram_reg_140__0_ ( .D(n6677), .CLK(clk), .Q(ram[2240]) );
  DFFPOSX1 ram_reg_139__15_ ( .D(n6676), .CLK(clk), .Q(ram[2239]) );
  DFFPOSX1 ram_reg_139__14_ ( .D(n6675), .CLK(clk), .Q(ram[2238]) );
  DFFPOSX1 ram_reg_139__13_ ( .D(n6674), .CLK(clk), .Q(ram[2237]) );
  DFFPOSX1 ram_reg_139__12_ ( .D(n6673), .CLK(clk), .Q(ram[2236]) );
  DFFPOSX1 ram_reg_139__11_ ( .D(n6672), .CLK(clk), .Q(ram[2235]) );
  DFFPOSX1 ram_reg_139__10_ ( .D(n6671), .CLK(clk), .Q(ram[2234]) );
  DFFPOSX1 ram_reg_139__9_ ( .D(n6670), .CLK(clk), .Q(ram[2233]) );
  DFFPOSX1 ram_reg_139__8_ ( .D(n6669), .CLK(clk), .Q(ram[2232]) );
  DFFPOSX1 ram_reg_139__7_ ( .D(n6668), .CLK(clk), .Q(ram[2231]) );
  DFFPOSX1 ram_reg_139__6_ ( .D(n6667), .CLK(clk), .Q(ram[2230]) );
  DFFPOSX1 ram_reg_139__5_ ( .D(n6666), .CLK(clk), .Q(ram[2229]) );
  DFFPOSX1 ram_reg_139__4_ ( .D(n6665), .CLK(clk), .Q(ram[2228]) );
  DFFPOSX1 ram_reg_139__3_ ( .D(n6664), .CLK(clk), .Q(ram[2227]) );
  DFFPOSX1 ram_reg_139__2_ ( .D(n6663), .CLK(clk), .Q(ram[2226]) );
  DFFPOSX1 ram_reg_139__1_ ( .D(n6662), .CLK(clk), .Q(ram[2225]) );
  DFFPOSX1 ram_reg_139__0_ ( .D(n6661), .CLK(clk), .Q(ram[2224]) );
  DFFPOSX1 ram_reg_138__15_ ( .D(n6660), .CLK(clk), .Q(ram[2223]) );
  DFFPOSX1 ram_reg_138__14_ ( .D(n6659), .CLK(clk), .Q(ram[2222]) );
  DFFPOSX1 ram_reg_138__13_ ( .D(n6658), .CLK(clk), .Q(ram[2221]) );
  DFFPOSX1 ram_reg_138__12_ ( .D(n6657), .CLK(clk), .Q(ram[2220]) );
  DFFPOSX1 ram_reg_138__11_ ( .D(n6656), .CLK(clk), .Q(ram[2219]) );
  DFFPOSX1 ram_reg_138__10_ ( .D(n6655), .CLK(clk), .Q(ram[2218]) );
  DFFPOSX1 ram_reg_138__9_ ( .D(n6654), .CLK(clk), .Q(ram[2217]) );
  DFFPOSX1 ram_reg_138__8_ ( .D(n6653), .CLK(clk), .Q(ram[2216]) );
  DFFPOSX1 ram_reg_138__7_ ( .D(n6652), .CLK(clk), .Q(ram[2215]) );
  DFFPOSX1 ram_reg_138__6_ ( .D(n6651), .CLK(clk), .Q(ram[2214]) );
  DFFPOSX1 ram_reg_138__5_ ( .D(n6650), .CLK(clk), .Q(ram[2213]) );
  DFFPOSX1 ram_reg_138__4_ ( .D(n6649), .CLK(clk), .Q(ram[2212]) );
  DFFPOSX1 ram_reg_138__3_ ( .D(n6648), .CLK(clk), .Q(ram[2211]) );
  DFFPOSX1 ram_reg_138__2_ ( .D(n6647), .CLK(clk), .Q(ram[2210]) );
  DFFPOSX1 ram_reg_138__1_ ( .D(n6646), .CLK(clk), .Q(ram[2209]) );
  DFFPOSX1 ram_reg_138__0_ ( .D(n6645), .CLK(clk), .Q(ram[2208]) );
  DFFPOSX1 ram_reg_137__15_ ( .D(n6644), .CLK(clk), .Q(ram[2207]) );
  DFFPOSX1 ram_reg_137__14_ ( .D(n6643), .CLK(clk), .Q(ram[2206]) );
  DFFPOSX1 ram_reg_137__13_ ( .D(n6642), .CLK(clk), .Q(ram[2205]) );
  DFFPOSX1 ram_reg_137__12_ ( .D(n6641), .CLK(clk), .Q(ram[2204]) );
  DFFPOSX1 ram_reg_137__11_ ( .D(n6640), .CLK(clk), .Q(ram[2203]) );
  DFFPOSX1 ram_reg_137__10_ ( .D(n6639), .CLK(clk), .Q(ram[2202]) );
  DFFPOSX1 ram_reg_137__9_ ( .D(n6638), .CLK(clk), .Q(ram[2201]) );
  DFFPOSX1 ram_reg_137__8_ ( .D(n6637), .CLK(clk), .Q(ram[2200]) );
  DFFPOSX1 ram_reg_137__7_ ( .D(n6636), .CLK(clk), .Q(ram[2199]) );
  DFFPOSX1 ram_reg_137__6_ ( .D(n6635), .CLK(clk), .Q(ram[2198]) );
  DFFPOSX1 ram_reg_137__5_ ( .D(n6634), .CLK(clk), .Q(ram[2197]) );
  DFFPOSX1 ram_reg_137__4_ ( .D(n6633), .CLK(clk), .Q(ram[2196]) );
  DFFPOSX1 ram_reg_137__3_ ( .D(n6632), .CLK(clk), .Q(ram[2195]) );
  DFFPOSX1 ram_reg_137__2_ ( .D(n6631), .CLK(clk), .Q(ram[2194]) );
  DFFPOSX1 ram_reg_137__1_ ( .D(n6630), .CLK(clk), .Q(ram[2193]) );
  DFFPOSX1 ram_reg_137__0_ ( .D(n6629), .CLK(clk), .Q(ram[2192]) );
  DFFPOSX1 ram_reg_136__15_ ( .D(n6628), .CLK(clk), .Q(ram[2191]) );
  DFFPOSX1 ram_reg_136__14_ ( .D(n6627), .CLK(clk), .Q(ram[2190]) );
  DFFPOSX1 ram_reg_136__13_ ( .D(n6626), .CLK(clk), .Q(ram[2189]) );
  DFFPOSX1 ram_reg_136__12_ ( .D(n6625), .CLK(clk), .Q(ram[2188]) );
  DFFPOSX1 ram_reg_136__11_ ( .D(n6624), .CLK(clk), .Q(ram[2187]) );
  DFFPOSX1 ram_reg_136__10_ ( .D(n6623), .CLK(clk), .Q(ram[2186]) );
  DFFPOSX1 ram_reg_136__9_ ( .D(n6622), .CLK(clk), .Q(ram[2185]) );
  DFFPOSX1 ram_reg_136__8_ ( .D(n6621), .CLK(clk), .Q(ram[2184]) );
  DFFPOSX1 ram_reg_136__7_ ( .D(n6620), .CLK(clk), .Q(ram[2183]) );
  DFFPOSX1 ram_reg_136__6_ ( .D(n6619), .CLK(clk), .Q(ram[2182]) );
  DFFPOSX1 ram_reg_136__5_ ( .D(n6618), .CLK(clk), .Q(ram[2181]) );
  DFFPOSX1 ram_reg_136__4_ ( .D(n6617), .CLK(clk), .Q(ram[2180]) );
  DFFPOSX1 ram_reg_136__3_ ( .D(n6616), .CLK(clk), .Q(ram[2179]) );
  DFFPOSX1 ram_reg_136__2_ ( .D(n6615), .CLK(clk), .Q(ram[2178]) );
  DFFPOSX1 ram_reg_136__1_ ( .D(n6614), .CLK(clk), .Q(ram[2177]) );
  DFFPOSX1 ram_reg_136__0_ ( .D(n6613), .CLK(clk), .Q(ram[2176]) );
  DFFPOSX1 ram_reg_135__15_ ( .D(n6612), .CLK(clk), .Q(ram[2175]) );
  DFFPOSX1 ram_reg_135__14_ ( .D(n6611), .CLK(clk), .Q(ram[2174]) );
  DFFPOSX1 ram_reg_135__13_ ( .D(n6610), .CLK(clk), .Q(ram[2173]) );
  DFFPOSX1 ram_reg_135__12_ ( .D(n6609), .CLK(clk), .Q(ram[2172]) );
  DFFPOSX1 ram_reg_135__11_ ( .D(n6608), .CLK(clk), .Q(ram[2171]) );
  DFFPOSX1 ram_reg_135__10_ ( .D(n6607), .CLK(clk), .Q(ram[2170]) );
  DFFPOSX1 ram_reg_135__9_ ( .D(n6606), .CLK(clk), .Q(ram[2169]) );
  DFFPOSX1 ram_reg_135__8_ ( .D(n6605), .CLK(clk), .Q(ram[2168]) );
  DFFPOSX1 ram_reg_135__7_ ( .D(n6604), .CLK(clk), .Q(ram[2167]) );
  DFFPOSX1 ram_reg_135__6_ ( .D(n6603), .CLK(clk), .Q(ram[2166]) );
  DFFPOSX1 ram_reg_135__5_ ( .D(n6602), .CLK(clk), .Q(ram[2165]) );
  DFFPOSX1 ram_reg_135__4_ ( .D(n6601), .CLK(clk), .Q(ram[2164]) );
  DFFPOSX1 ram_reg_135__3_ ( .D(n6600), .CLK(clk), .Q(ram[2163]) );
  DFFPOSX1 ram_reg_135__2_ ( .D(n6599), .CLK(clk), .Q(ram[2162]) );
  DFFPOSX1 ram_reg_135__1_ ( .D(n6598), .CLK(clk), .Q(ram[2161]) );
  DFFPOSX1 ram_reg_135__0_ ( .D(n6597), .CLK(clk), .Q(ram[2160]) );
  DFFPOSX1 ram_reg_134__15_ ( .D(n6596), .CLK(clk), .Q(ram[2159]) );
  DFFPOSX1 ram_reg_134__14_ ( .D(n6595), .CLK(clk), .Q(ram[2158]) );
  DFFPOSX1 ram_reg_134__13_ ( .D(n6594), .CLK(clk), .Q(ram[2157]) );
  DFFPOSX1 ram_reg_134__12_ ( .D(n6593), .CLK(clk), .Q(ram[2156]) );
  DFFPOSX1 ram_reg_134__11_ ( .D(n6592), .CLK(clk), .Q(ram[2155]) );
  DFFPOSX1 ram_reg_134__10_ ( .D(n6591), .CLK(clk), .Q(ram[2154]) );
  DFFPOSX1 ram_reg_134__9_ ( .D(n6590), .CLK(clk), .Q(ram[2153]) );
  DFFPOSX1 ram_reg_134__8_ ( .D(n6589), .CLK(clk), .Q(ram[2152]) );
  DFFPOSX1 ram_reg_134__7_ ( .D(n6588), .CLK(clk), .Q(ram[2151]) );
  DFFPOSX1 ram_reg_134__6_ ( .D(n6587), .CLK(clk), .Q(ram[2150]) );
  DFFPOSX1 ram_reg_134__5_ ( .D(n6586), .CLK(clk), .Q(ram[2149]) );
  DFFPOSX1 ram_reg_134__4_ ( .D(n6585), .CLK(clk), .Q(ram[2148]) );
  DFFPOSX1 ram_reg_134__3_ ( .D(n6584), .CLK(clk), .Q(ram[2147]) );
  DFFPOSX1 ram_reg_134__2_ ( .D(n6583), .CLK(clk), .Q(ram[2146]) );
  DFFPOSX1 ram_reg_134__1_ ( .D(n6582), .CLK(clk), .Q(ram[2145]) );
  DFFPOSX1 ram_reg_134__0_ ( .D(n6581), .CLK(clk), .Q(ram[2144]) );
  DFFPOSX1 ram_reg_133__15_ ( .D(n6580), .CLK(clk), .Q(ram[2143]) );
  DFFPOSX1 ram_reg_133__14_ ( .D(n6579), .CLK(clk), .Q(ram[2142]) );
  DFFPOSX1 ram_reg_133__13_ ( .D(n6578), .CLK(clk), .Q(ram[2141]) );
  DFFPOSX1 ram_reg_133__12_ ( .D(n6577), .CLK(clk), .Q(ram[2140]) );
  DFFPOSX1 ram_reg_133__11_ ( .D(n6576), .CLK(clk), .Q(ram[2139]) );
  DFFPOSX1 ram_reg_133__10_ ( .D(n6575), .CLK(clk), .Q(ram[2138]) );
  DFFPOSX1 ram_reg_133__9_ ( .D(n6574), .CLK(clk), .Q(ram[2137]) );
  DFFPOSX1 ram_reg_133__8_ ( .D(n6573), .CLK(clk), .Q(ram[2136]) );
  DFFPOSX1 ram_reg_133__7_ ( .D(n6572), .CLK(clk), .Q(ram[2135]) );
  DFFPOSX1 ram_reg_133__6_ ( .D(n6571), .CLK(clk), .Q(ram[2134]) );
  DFFPOSX1 ram_reg_133__5_ ( .D(n6570), .CLK(clk), .Q(ram[2133]) );
  DFFPOSX1 ram_reg_133__4_ ( .D(n6569), .CLK(clk), .Q(ram[2132]) );
  DFFPOSX1 ram_reg_133__3_ ( .D(n6568), .CLK(clk), .Q(ram[2131]) );
  DFFPOSX1 ram_reg_133__2_ ( .D(n6567), .CLK(clk), .Q(ram[2130]) );
  DFFPOSX1 ram_reg_133__1_ ( .D(n6566), .CLK(clk), .Q(ram[2129]) );
  DFFPOSX1 ram_reg_133__0_ ( .D(n6565), .CLK(clk), .Q(ram[2128]) );
  DFFPOSX1 ram_reg_132__15_ ( .D(n6564), .CLK(clk), .Q(ram[2127]) );
  DFFPOSX1 ram_reg_132__14_ ( .D(n6563), .CLK(clk), .Q(ram[2126]) );
  DFFPOSX1 ram_reg_132__13_ ( .D(n6562), .CLK(clk), .Q(ram[2125]) );
  DFFPOSX1 ram_reg_132__12_ ( .D(n6561), .CLK(clk), .Q(ram[2124]) );
  DFFPOSX1 ram_reg_132__11_ ( .D(n6560), .CLK(clk), .Q(ram[2123]) );
  DFFPOSX1 ram_reg_132__10_ ( .D(n6559), .CLK(clk), .Q(ram[2122]) );
  DFFPOSX1 ram_reg_132__9_ ( .D(n6558), .CLK(clk), .Q(ram[2121]) );
  DFFPOSX1 ram_reg_132__8_ ( .D(n6557), .CLK(clk), .Q(ram[2120]) );
  DFFPOSX1 ram_reg_132__7_ ( .D(n6556), .CLK(clk), .Q(ram[2119]) );
  DFFPOSX1 ram_reg_132__6_ ( .D(n6555), .CLK(clk), .Q(ram[2118]) );
  DFFPOSX1 ram_reg_132__5_ ( .D(n6554), .CLK(clk), .Q(ram[2117]) );
  DFFPOSX1 ram_reg_132__4_ ( .D(n6553), .CLK(clk), .Q(ram[2116]) );
  DFFPOSX1 ram_reg_132__3_ ( .D(n6552), .CLK(clk), .Q(ram[2115]) );
  DFFPOSX1 ram_reg_132__2_ ( .D(n6551), .CLK(clk), .Q(ram[2114]) );
  DFFPOSX1 ram_reg_132__1_ ( .D(n6550), .CLK(clk), .Q(ram[2113]) );
  DFFPOSX1 ram_reg_132__0_ ( .D(n6549), .CLK(clk), .Q(ram[2112]) );
  DFFPOSX1 ram_reg_131__15_ ( .D(n6548), .CLK(clk), .Q(ram[2111]) );
  DFFPOSX1 ram_reg_131__14_ ( .D(n6547), .CLK(clk), .Q(ram[2110]) );
  DFFPOSX1 ram_reg_131__13_ ( .D(n6546), .CLK(clk), .Q(ram[2109]) );
  DFFPOSX1 ram_reg_131__12_ ( .D(n6545), .CLK(clk), .Q(ram[2108]) );
  DFFPOSX1 ram_reg_131__11_ ( .D(n6544), .CLK(clk), .Q(ram[2107]) );
  DFFPOSX1 ram_reg_131__10_ ( .D(n6543), .CLK(clk), .Q(ram[2106]) );
  DFFPOSX1 ram_reg_131__9_ ( .D(n6542), .CLK(clk), .Q(ram[2105]) );
  DFFPOSX1 ram_reg_131__8_ ( .D(n6541), .CLK(clk), .Q(ram[2104]) );
  DFFPOSX1 ram_reg_131__7_ ( .D(n6540), .CLK(clk), .Q(ram[2103]) );
  DFFPOSX1 ram_reg_131__6_ ( .D(n6539), .CLK(clk), .Q(ram[2102]) );
  DFFPOSX1 ram_reg_131__5_ ( .D(n6538), .CLK(clk), .Q(ram[2101]) );
  DFFPOSX1 ram_reg_131__4_ ( .D(n6537), .CLK(clk), .Q(ram[2100]) );
  DFFPOSX1 ram_reg_131__3_ ( .D(n6536), .CLK(clk), .Q(ram[2099]) );
  DFFPOSX1 ram_reg_131__2_ ( .D(n6535), .CLK(clk), .Q(ram[2098]) );
  DFFPOSX1 ram_reg_131__1_ ( .D(n6534), .CLK(clk), .Q(ram[2097]) );
  DFFPOSX1 ram_reg_131__0_ ( .D(n6533), .CLK(clk), .Q(ram[2096]) );
  DFFPOSX1 ram_reg_130__15_ ( .D(n6532), .CLK(clk), .Q(ram[2095]) );
  DFFPOSX1 ram_reg_130__14_ ( .D(n6531), .CLK(clk), .Q(ram[2094]) );
  DFFPOSX1 ram_reg_130__13_ ( .D(n6530), .CLK(clk), .Q(ram[2093]) );
  DFFPOSX1 ram_reg_130__12_ ( .D(n6529), .CLK(clk), .Q(ram[2092]) );
  DFFPOSX1 ram_reg_130__11_ ( .D(n6528), .CLK(clk), .Q(ram[2091]) );
  DFFPOSX1 ram_reg_130__10_ ( .D(n6527), .CLK(clk), .Q(ram[2090]) );
  DFFPOSX1 ram_reg_130__9_ ( .D(n6526), .CLK(clk), .Q(ram[2089]) );
  DFFPOSX1 ram_reg_130__8_ ( .D(n6525), .CLK(clk), .Q(ram[2088]) );
  DFFPOSX1 ram_reg_130__7_ ( .D(n6524), .CLK(clk), .Q(ram[2087]) );
  DFFPOSX1 ram_reg_130__6_ ( .D(n6523), .CLK(clk), .Q(ram[2086]) );
  DFFPOSX1 ram_reg_130__5_ ( .D(n6522), .CLK(clk), .Q(ram[2085]) );
  DFFPOSX1 ram_reg_130__4_ ( .D(n6521), .CLK(clk), .Q(ram[2084]) );
  DFFPOSX1 ram_reg_130__3_ ( .D(n6520), .CLK(clk), .Q(ram[2083]) );
  DFFPOSX1 ram_reg_130__2_ ( .D(n6519), .CLK(clk), .Q(ram[2082]) );
  DFFPOSX1 ram_reg_130__1_ ( .D(n6518), .CLK(clk), .Q(ram[2081]) );
  DFFPOSX1 ram_reg_130__0_ ( .D(n6517), .CLK(clk), .Q(ram[2080]) );
  DFFPOSX1 ram_reg_129__15_ ( .D(n6516), .CLK(clk), .Q(ram[2079]) );
  DFFPOSX1 ram_reg_129__14_ ( .D(n6515), .CLK(clk), .Q(ram[2078]) );
  DFFPOSX1 ram_reg_129__13_ ( .D(n6514), .CLK(clk), .Q(ram[2077]) );
  DFFPOSX1 ram_reg_129__12_ ( .D(n6513), .CLK(clk), .Q(ram[2076]) );
  DFFPOSX1 ram_reg_129__11_ ( .D(n6512), .CLK(clk), .Q(ram[2075]) );
  DFFPOSX1 ram_reg_129__10_ ( .D(n6511), .CLK(clk), .Q(ram[2074]) );
  DFFPOSX1 ram_reg_129__9_ ( .D(n6510), .CLK(clk), .Q(ram[2073]) );
  DFFPOSX1 ram_reg_129__8_ ( .D(n6509), .CLK(clk), .Q(ram[2072]) );
  DFFPOSX1 ram_reg_129__7_ ( .D(n6508), .CLK(clk), .Q(ram[2071]) );
  DFFPOSX1 ram_reg_129__6_ ( .D(n6507), .CLK(clk), .Q(ram[2070]) );
  DFFPOSX1 ram_reg_129__5_ ( .D(n6506), .CLK(clk), .Q(ram[2069]) );
  DFFPOSX1 ram_reg_129__4_ ( .D(n6505), .CLK(clk), .Q(ram[2068]) );
  DFFPOSX1 ram_reg_129__3_ ( .D(n6504), .CLK(clk), .Q(ram[2067]) );
  DFFPOSX1 ram_reg_129__2_ ( .D(n6503), .CLK(clk), .Q(ram[2066]) );
  DFFPOSX1 ram_reg_129__1_ ( .D(n6502), .CLK(clk), .Q(ram[2065]) );
  DFFPOSX1 ram_reg_129__0_ ( .D(n6501), .CLK(clk), .Q(ram[2064]) );
  DFFPOSX1 ram_reg_128__15_ ( .D(n6500), .CLK(clk), .Q(ram[2063]) );
  DFFPOSX1 ram_reg_128__14_ ( .D(n6499), .CLK(clk), .Q(ram[2062]) );
  DFFPOSX1 ram_reg_128__13_ ( .D(n6498), .CLK(clk), .Q(ram[2061]) );
  DFFPOSX1 ram_reg_128__12_ ( .D(n6497), .CLK(clk), .Q(ram[2060]) );
  DFFPOSX1 ram_reg_128__11_ ( .D(n6496), .CLK(clk), .Q(ram[2059]) );
  DFFPOSX1 ram_reg_128__10_ ( .D(n6495), .CLK(clk), .Q(ram[2058]) );
  DFFPOSX1 ram_reg_128__9_ ( .D(n6494), .CLK(clk), .Q(ram[2057]) );
  DFFPOSX1 ram_reg_128__8_ ( .D(n6493), .CLK(clk), .Q(ram[2056]) );
  DFFPOSX1 ram_reg_128__7_ ( .D(n6492), .CLK(clk), .Q(ram[2055]) );
  DFFPOSX1 ram_reg_128__6_ ( .D(n6491), .CLK(clk), .Q(ram[2054]) );
  DFFPOSX1 ram_reg_128__5_ ( .D(n6490), .CLK(clk), .Q(ram[2053]) );
  DFFPOSX1 ram_reg_128__4_ ( .D(n6489), .CLK(clk), .Q(ram[2052]) );
  DFFPOSX1 ram_reg_128__3_ ( .D(n6488), .CLK(clk), .Q(ram[2051]) );
  DFFPOSX1 ram_reg_128__2_ ( .D(n6487), .CLK(clk), .Q(ram[2050]) );
  DFFPOSX1 ram_reg_128__1_ ( .D(n6486), .CLK(clk), .Q(ram[2049]) );
  DFFPOSX1 ram_reg_128__0_ ( .D(n6485), .CLK(clk), .Q(ram[2048]) );
  DFFPOSX1 ram_reg_127__15_ ( .D(n6484), .CLK(clk), .Q(ram[2047]) );
  DFFPOSX1 ram_reg_127__14_ ( .D(n6483), .CLK(clk), .Q(ram[2046]) );
  DFFPOSX1 ram_reg_127__13_ ( .D(n6482), .CLK(clk), .Q(ram[2045]) );
  DFFPOSX1 ram_reg_127__12_ ( .D(n6481), .CLK(clk), .Q(ram[2044]) );
  DFFPOSX1 ram_reg_127__11_ ( .D(n6480), .CLK(clk), .Q(ram[2043]) );
  DFFPOSX1 ram_reg_127__10_ ( .D(n6479), .CLK(clk), .Q(ram[2042]) );
  DFFPOSX1 ram_reg_127__9_ ( .D(n6478), .CLK(clk), .Q(ram[2041]) );
  DFFPOSX1 ram_reg_127__8_ ( .D(n6477), .CLK(clk), .Q(ram[2040]) );
  DFFPOSX1 ram_reg_127__7_ ( .D(n6476), .CLK(clk), .Q(ram[2039]) );
  DFFPOSX1 ram_reg_127__6_ ( .D(n6475), .CLK(clk), .Q(ram[2038]) );
  DFFPOSX1 ram_reg_127__5_ ( .D(n6474), .CLK(clk), .Q(ram[2037]) );
  DFFPOSX1 ram_reg_127__4_ ( .D(n6473), .CLK(clk), .Q(ram[2036]) );
  DFFPOSX1 ram_reg_127__3_ ( .D(n6472), .CLK(clk), .Q(ram[2035]) );
  DFFPOSX1 ram_reg_127__2_ ( .D(n6471), .CLK(clk), .Q(ram[2034]) );
  DFFPOSX1 ram_reg_127__1_ ( .D(n6470), .CLK(clk), .Q(ram[2033]) );
  DFFPOSX1 ram_reg_127__0_ ( .D(n6469), .CLK(clk), .Q(ram[2032]) );
  DFFPOSX1 ram_reg_126__15_ ( .D(n6468), .CLK(clk), .Q(ram[2031]) );
  DFFPOSX1 ram_reg_126__14_ ( .D(n6467), .CLK(clk), .Q(ram[2030]) );
  DFFPOSX1 ram_reg_126__13_ ( .D(n6466), .CLK(clk), .Q(ram[2029]) );
  DFFPOSX1 ram_reg_126__12_ ( .D(n6465), .CLK(clk), .Q(ram[2028]) );
  DFFPOSX1 ram_reg_126__11_ ( .D(n6464), .CLK(clk), .Q(ram[2027]) );
  DFFPOSX1 ram_reg_126__10_ ( .D(n6463), .CLK(clk), .Q(ram[2026]) );
  DFFPOSX1 ram_reg_126__9_ ( .D(n6462), .CLK(clk), .Q(ram[2025]) );
  DFFPOSX1 ram_reg_126__8_ ( .D(n6461), .CLK(clk), .Q(ram[2024]) );
  DFFPOSX1 ram_reg_126__7_ ( .D(n6460), .CLK(clk), .Q(ram[2023]) );
  DFFPOSX1 ram_reg_126__6_ ( .D(n6459), .CLK(clk), .Q(ram[2022]) );
  DFFPOSX1 ram_reg_126__5_ ( .D(n6458), .CLK(clk), .Q(ram[2021]) );
  DFFPOSX1 ram_reg_126__4_ ( .D(n6457), .CLK(clk), .Q(ram[2020]) );
  DFFPOSX1 ram_reg_126__3_ ( .D(n6456), .CLK(clk), .Q(ram[2019]) );
  DFFPOSX1 ram_reg_126__2_ ( .D(n6455), .CLK(clk), .Q(ram[2018]) );
  DFFPOSX1 ram_reg_126__1_ ( .D(n6454), .CLK(clk), .Q(ram[2017]) );
  DFFPOSX1 ram_reg_126__0_ ( .D(n6453), .CLK(clk), .Q(ram[2016]) );
  DFFPOSX1 ram_reg_125__15_ ( .D(n6452), .CLK(clk), .Q(ram[2015]) );
  DFFPOSX1 ram_reg_125__14_ ( .D(n6451), .CLK(clk), .Q(ram[2014]) );
  DFFPOSX1 ram_reg_125__13_ ( .D(n6450), .CLK(clk), .Q(ram[2013]) );
  DFFPOSX1 ram_reg_125__12_ ( .D(n6449), .CLK(clk), .Q(ram[2012]) );
  DFFPOSX1 ram_reg_125__11_ ( .D(n6448), .CLK(clk), .Q(ram[2011]) );
  DFFPOSX1 ram_reg_125__10_ ( .D(n6447), .CLK(clk), .Q(ram[2010]) );
  DFFPOSX1 ram_reg_125__9_ ( .D(n6446), .CLK(clk), .Q(ram[2009]) );
  DFFPOSX1 ram_reg_125__8_ ( .D(n6445), .CLK(clk), .Q(ram[2008]) );
  DFFPOSX1 ram_reg_125__7_ ( .D(n6444), .CLK(clk), .Q(ram[2007]) );
  DFFPOSX1 ram_reg_125__6_ ( .D(n6443), .CLK(clk), .Q(ram[2006]) );
  DFFPOSX1 ram_reg_125__5_ ( .D(n6442), .CLK(clk), .Q(ram[2005]) );
  DFFPOSX1 ram_reg_125__4_ ( .D(n6441), .CLK(clk), .Q(ram[2004]) );
  DFFPOSX1 ram_reg_125__3_ ( .D(n6440), .CLK(clk), .Q(ram[2003]) );
  DFFPOSX1 ram_reg_125__2_ ( .D(n6439), .CLK(clk), .Q(ram[2002]) );
  DFFPOSX1 ram_reg_125__1_ ( .D(n6438), .CLK(clk), .Q(ram[2001]) );
  DFFPOSX1 ram_reg_125__0_ ( .D(n6437), .CLK(clk), .Q(ram[2000]) );
  DFFPOSX1 ram_reg_124__15_ ( .D(n6436), .CLK(clk), .Q(ram[1999]) );
  DFFPOSX1 ram_reg_124__14_ ( .D(n6435), .CLK(clk), .Q(ram[1998]) );
  DFFPOSX1 ram_reg_124__13_ ( .D(n6434), .CLK(clk), .Q(ram[1997]) );
  DFFPOSX1 ram_reg_124__12_ ( .D(n6433), .CLK(clk), .Q(ram[1996]) );
  DFFPOSX1 ram_reg_124__11_ ( .D(n6432), .CLK(clk), .Q(ram[1995]) );
  DFFPOSX1 ram_reg_124__10_ ( .D(n6431), .CLK(clk), .Q(ram[1994]) );
  DFFPOSX1 ram_reg_124__9_ ( .D(n6430), .CLK(clk), .Q(ram[1993]) );
  DFFPOSX1 ram_reg_124__8_ ( .D(n6429), .CLK(clk), .Q(ram[1992]) );
  DFFPOSX1 ram_reg_124__7_ ( .D(n6428), .CLK(clk), .Q(ram[1991]) );
  DFFPOSX1 ram_reg_124__6_ ( .D(n6427), .CLK(clk), .Q(ram[1990]) );
  DFFPOSX1 ram_reg_124__5_ ( .D(n6426), .CLK(clk), .Q(ram[1989]) );
  DFFPOSX1 ram_reg_124__4_ ( .D(n6425), .CLK(clk), .Q(ram[1988]) );
  DFFPOSX1 ram_reg_124__3_ ( .D(n6424), .CLK(clk), .Q(ram[1987]) );
  DFFPOSX1 ram_reg_124__2_ ( .D(n6423), .CLK(clk), .Q(ram[1986]) );
  DFFPOSX1 ram_reg_124__1_ ( .D(n6422), .CLK(clk), .Q(ram[1985]) );
  DFFPOSX1 ram_reg_124__0_ ( .D(n6421), .CLK(clk), .Q(ram[1984]) );
  DFFPOSX1 ram_reg_123__15_ ( .D(n6420), .CLK(clk), .Q(ram[1983]) );
  DFFPOSX1 ram_reg_123__14_ ( .D(n6419), .CLK(clk), .Q(ram[1982]) );
  DFFPOSX1 ram_reg_123__13_ ( .D(n6418), .CLK(clk), .Q(ram[1981]) );
  DFFPOSX1 ram_reg_123__12_ ( .D(n6417), .CLK(clk), .Q(ram[1980]) );
  DFFPOSX1 ram_reg_123__11_ ( .D(n6416), .CLK(clk), .Q(ram[1979]) );
  DFFPOSX1 ram_reg_123__10_ ( .D(n6415), .CLK(clk), .Q(ram[1978]) );
  DFFPOSX1 ram_reg_123__9_ ( .D(n6414), .CLK(clk), .Q(ram[1977]) );
  DFFPOSX1 ram_reg_123__8_ ( .D(n6413), .CLK(clk), .Q(ram[1976]) );
  DFFPOSX1 ram_reg_123__7_ ( .D(n6412), .CLK(clk), .Q(ram[1975]) );
  DFFPOSX1 ram_reg_123__6_ ( .D(n6411), .CLK(clk), .Q(ram[1974]) );
  DFFPOSX1 ram_reg_123__5_ ( .D(n6410), .CLK(clk), .Q(ram[1973]) );
  DFFPOSX1 ram_reg_123__4_ ( .D(n6409), .CLK(clk), .Q(ram[1972]) );
  DFFPOSX1 ram_reg_123__3_ ( .D(n6408), .CLK(clk), .Q(ram[1971]) );
  DFFPOSX1 ram_reg_123__2_ ( .D(n6407), .CLK(clk), .Q(ram[1970]) );
  DFFPOSX1 ram_reg_123__1_ ( .D(n6406), .CLK(clk), .Q(ram[1969]) );
  DFFPOSX1 ram_reg_123__0_ ( .D(n6405), .CLK(clk), .Q(ram[1968]) );
  DFFPOSX1 ram_reg_122__15_ ( .D(n6404), .CLK(clk), .Q(ram[1967]) );
  DFFPOSX1 ram_reg_122__14_ ( .D(n6403), .CLK(clk), .Q(ram[1966]) );
  DFFPOSX1 ram_reg_122__13_ ( .D(n6402), .CLK(clk), .Q(ram[1965]) );
  DFFPOSX1 ram_reg_122__12_ ( .D(n6401), .CLK(clk), .Q(ram[1964]) );
  DFFPOSX1 ram_reg_122__11_ ( .D(n6400), .CLK(clk), .Q(ram[1963]) );
  DFFPOSX1 ram_reg_122__10_ ( .D(n6399), .CLK(clk), .Q(ram[1962]) );
  DFFPOSX1 ram_reg_122__9_ ( .D(n6398), .CLK(clk), .Q(ram[1961]) );
  DFFPOSX1 ram_reg_122__8_ ( .D(n6397), .CLK(clk), .Q(ram[1960]) );
  DFFPOSX1 ram_reg_122__7_ ( .D(n6396), .CLK(clk), .Q(ram[1959]) );
  DFFPOSX1 ram_reg_122__6_ ( .D(n6395), .CLK(clk), .Q(ram[1958]) );
  DFFPOSX1 ram_reg_122__5_ ( .D(n6394), .CLK(clk), .Q(ram[1957]) );
  DFFPOSX1 ram_reg_122__4_ ( .D(n6393), .CLK(clk), .Q(ram[1956]) );
  DFFPOSX1 ram_reg_122__3_ ( .D(n6392), .CLK(clk), .Q(ram[1955]) );
  DFFPOSX1 ram_reg_122__2_ ( .D(n6391), .CLK(clk), .Q(ram[1954]) );
  DFFPOSX1 ram_reg_122__1_ ( .D(n6390), .CLK(clk), .Q(ram[1953]) );
  DFFPOSX1 ram_reg_122__0_ ( .D(n6389), .CLK(clk), .Q(ram[1952]) );
  DFFPOSX1 ram_reg_121__15_ ( .D(n6388), .CLK(clk), .Q(ram[1951]) );
  DFFPOSX1 ram_reg_121__14_ ( .D(n6387), .CLK(clk), .Q(ram[1950]) );
  DFFPOSX1 ram_reg_121__13_ ( .D(n6386), .CLK(clk), .Q(ram[1949]) );
  DFFPOSX1 ram_reg_121__12_ ( .D(n6385), .CLK(clk), .Q(ram[1948]) );
  DFFPOSX1 ram_reg_121__11_ ( .D(n6384), .CLK(clk), .Q(ram[1947]) );
  DFFPOSX1 ram_reg_121__10_ ( .D(n6383), .CLK(clk), .Q(ram[1946]) );
  DFFPOSX1 ram_reg_121__9_ ( .D(n6382), .CLK(clk), .Q(ram[1945]) );
  DFFPOSX1 ram_reg_121__8_ ( .D(n6381), .CLK(clk), .Q(ram[1944]) );
  DFFPOSX1 ram_reg_121__7_ ( .D(n6380), .CLK(clk), .Q(ram[1943]) );
  DFFPOSX1 ram_reg_121__6_ ( .D(n6379), .CLK(clk), .Q(ram[1942]) );
  DFFPOSX1 ram_reg_121__5_ ( .D(n6378), .CLK(clk), .Q(ram[1941]) );
  DFFPOSX1 ram_reg_121__4_ ( .D(n6377), .CLK(clk), .Q(ram[1940]) );
  DFFPOSX1 ram_reg_121__3_ ( .D(n6376), .CLK(clk), .Q(ram[1939]) );
  DFFPOSX1 ram_reg_121__2_ ( .D(n6375), .CLK(clk), .Q(ram[1938]) );
  DFFPOSX1 ram_reg_121__1_ ( .D(n6374), .CLK(clk), .Q(ram[1937]) );
  DFFPOSX1 ram_reg_121__0_ ( .D(n6373), .CLK(clk), .Q(ram[1936]) );
  DFFPOSX1 ram_reg_120__15_ ( .D(n6372), .CLK(clk), .Q(ram[1935]) );
  DFFPOSX1 ram_reg_120__14_ ( .D(n6371), .CLK(clk), .Q(ram[1934]) );
  DFFPOSX1 ram_reg_120__13_ ( .D(n6370), .CLK(clk), .Q(ram[1933]) );
  DFFPOSX1 ram_reg_120__12_ ( .D(n6369), .CLK(clk), .Q(ram[1932]) );
  DFFPOSX1 ram_reg_120__11_ ( .D(n6368), .CLK(clk), .Q(ram[1931]) );
  DFFPOSX1 ram_reg_120__10_ ( .D(n6367), .CLK(clk), .Q(ram[1930]) );
  DFFPOSX1 ram_reg_120__9_ ( .D(n6366), .CLK(clk), .Q(ram[1929]) );
  DFFPOSX1 ram_reg_120__8_ ( .D(n6365), .CLK(clk), .Q(ram[1928]) );
  DFFPOSX1 ram_reg_120__7_ ( .D(n6364), .CLK(clk), .Q(ram[1927]) );
  DFFPOSX1 ram_reg_120__6_ ( .D(n6363), .CLK(clk), .Q(ram[1926]) );
  DFFPOSX1 ram_reg_120__5_ ( .D(n6362), .CLK(clk), .Q(ram[1925]) );
  DFFPOSX1 ram_reg_120__4_ ( .D(n6361), .CLK(clk), .Q(ram[1924]) );
  DFFPOSX1 ram_reg_120__3_ ( .D(n6360), .CLK(clk), .Q(ram[1923]) );
  DFFPOSX1 ram_reg_120__2_ ( .D(n6359), .CLK(clk), .Q(ram[1922]) );
  DFFPOSX1 ram_reg_120__1_ ( .D(n6358), .CLK(clk), .Q(ram[1921]) );
  DFFPOSX1 ram_reg_120__0_ ( .D(n6357), .CLK(clk), .Q(ram[1920]) );
  DFFPOSX1 ram_reg_119__15_ ( .D(n6356), .CLK(clk), .Q(ram[1919]) );
  DFFPOSX1 ram_reg_119__14_ ( .D(n6355), .CLK(clk), .Q(ram[1918]) );
  DFFPOSX1 ram_reg_119__13_ ( .D(n6354), .CLK(clk), .Q(ram[1917]) );
  DFFPOSX1 ram_reg_119__12_ ( .D(n6353), .CLK(clk), .Q(ram[1916]) );
  DFFPOSX1 ram_reg_119__11_ ( .D(n6352), .CLK(clk), .Q(ram[1915]) );
  DFFPOSX1 ram_reg_119__10_ ( .D(n6351), .CLK(clk), .Q(ram[1914]) );
  DFFPOSX1 ram_reg_119__9_ ( .D(n6350), .CLK(clk), .Q(ram[1913]) );
  DFFPOSX1 ram_reg_119__8_ ( .D(n6349), .CLK(clk), .Q(ram[1912]) );
  DFFPOSX1 ram_reg_119__7_ ( .D(n6348), .CLK(clk), .Q(ram[1911]) );
  DFFPOSX1 ram_reg_119__6_ ( .D(n6347), .CLK(clk), .Q(ram[1910]) );
  DFFPOSX1 ram_reg_119__5_ ( .D(n6346), .CLK(clk), .Q(ram[1909]) );
  DFFPOSX1 ram_reg_119__4_ ( .D(n6345), .CLK(clk), .Q(ram[1908]) );
  DFFPOSX1 ram_reg_119__3_ ( .D(n6344), .CLK(clk), .Q(ram[1907]) );
  DFFPOSX1 ram_reg_119__2_ ( .D(n6343), .CLK(clk), .Q(ram[1906]) );
  DFFPOSX1 ram_reg_119__1_ ( .D(n6342), .CLK(clk), .Q(ram[1905]) );
  DFFPOSX1 ram_reg_119__0_ ( .D(n6341), .CLK(clk), .Q(ram[1904]) );
  DFFPOSX1 ram_reg_118__15_ ( .D(n6340), .CLK(clk), .Q(ram[1903]) );
  DFFPOSX1 ram_reg_118__14_ ( .D(n6339), .CLK(clk), .Q(ram[1902]) );
  DFFPOSX1 ram_reg_118__13_ ( .D(n6338), .CLK(clk), .Q(ram[1901]) );
  DFFPOSX1 ram_reg_118__12_ ( .D(n6337), .CLK(clk), .Q(ram[1900]) );
  DFFPOSX1 ram_reg_118__11_ ( .D(n6336), .CLK(clk), .Q(ram[1899]) );
  DFFPOSX1 ram_reg_118__10_ ( .D(n6335), .CLK(clk), .Q(ram[1898]) );
  DFFPOSX1 ram_reg_118__9_ ( .D(n6334), .CLK(clk), .Q(ram[1897]) );
  DFFPOSX1 ram_reg_118__8_ ( .D(n6333), .CLK(clk), .Q(ram[1896]) );
  DFFPOSX1 ram_reg_118__7_ ( .D(n6332), .CLK(clk), .Q(ram[1895]) );
  DFFPOSX1 ram_reg_118__6_ ( .D(n6331), .CLK(clk), .Q(ram[1894]) );
  DFFPOSX1 ram_reg_118__5_ ( .D(n6330), .CLK(clk), .Q(ram[1893]) );
  DFFPOSX1 ram_reg_118__4_ ( .D(n6329), .CLK(clk), .Q(ram[1892]) );
  DFFPOSX1 ram_reg_118__3_ ( .D(n6328), .CLK(clk), .Q(ram[1891]) );
  DFFPOSX1 ram_reg_118__2_ ( .D(n6327), .CLK(clk), .Q(ram[1890]) );
  DFFPOSX1 ram_reg_118__1_ ( .D(n6326), .CLK(clk), .Q(ram[1889]) );
  DFFPOSX1 ram_reg_118__0_ ( .D(n6325), .CLK(clk), .Q(ram[1888]) );
  DFFPOSX1 ram_reg_117__15_ ( .D(n6324), .CLK(clk), .Q(ram[1887]) );
  DFFPOSX1 ram_reg_117__14_ ( .D(n6323), .CLK(clk), .Q(ram[1886]) );
  DFFPOSX1 ram_reg_117__13_ ( .D(n6322), .CLK(clk), .Q(ram[1885]) );
  DFFPOSX1 ram_reg_117__12_ ( .D(n6321), .CLK(clk), .Q(ram[1884]) );
  DFFPOSX1 ram_reg_117__11_ ( .D(n6320), .CLK(clk), .Q(ram[1883]) );
  DFFPOSX1 ram_reg_117__10_ ( .D(n6319), .CLK(clk), .Q(ram[1882]) );
  DFFPOSX1 ram_reg_117__9_ ( .D(n6318), .CLK(clk), .Q(ram[1881]) );
  DFFPOSX1 ram_reg_117__8_ ( .D(n6317), .CLK(clk), .Q(ram[1880]) );
  DFFPOSX1 ram_reg_117__7_ ( .D(n6316), .CLK(clk), .Q(ram[1879]) );
  DFFPOSX1 ram_reg_117__6_ ( .D(n6315), .CLK(clk), .Q(ram[1878]) );
  DFFPOSX1 ram_reg_117__5_ ( .D(n6314), .CLK(clk), .Q(ram[1877]) );
  DFFPOSX1 ram_reg_117__4_ ( .D(n6313), .CLK(clk), .Q(ram[1876]) );
  DFFPOSX1 ram_reg_117__3_ ( .D(n6312), .CLK(clk), .Q(ram[1875]) );
  DFFPOSX1 ram_reg_117__2_ ( .D(n6311), .CLK(clk), .Q(ram[1874]) );
  DFFPOSX1 ram_reg_117__1_ ( .D(n6310), .CLK(clk), .Q(ram[1873]) );
  DFFPOSX1 ram_reg_117__0_ ( .D(n6309), .CLK(clk), .Q(ram[1872]) );
  DFFPOSX1 ram_reg_116__15_ ( .D(n6308), .CLK(clk), .Q(ram[1871]) );
  DFFPOSX1 ram_reg_116__14_ ( .D(n6307), .CLK(clk), .Q(ram[1870]) );
  DFFPOSX1 ram_reg_116__13_ ( .D(n6306), .CLK(clk), .Q(ram[1869]) );
  DFFPOSX1 ram_reg_116__12_ ( .D(n6305), .CLK(clk), .Q(ram[1868]) );
  DFFPOSX1 ram_reg_116__11_ ( .D(n6304), .CLK(clk), .Q(ram[1867]) );
  DFFPOSX1 ram_reg_116__10_ ( .D(n6303), .CLK(clk), .Q(ram[1866]) );
  DFFPOSX1 ram_reg_116__9_ ( .D(n6302), .CLK(clk), .Q(ram[1865]) );
  DFFPOSX1 ram_reg_116__8_ ( .D(n6301), .CLK(clk), .Q(ram[1864]) );
  DFFPOSX1 ram_reg_116__7_ ( .D(n6300), .CLK(clk), .Q(ram[1863]) );
  DFFPOSX1 ram_reg_116__6_ ( .D(n6299), .CLK(clk), .Q(ram[1862]) );
  DFFPOSX1 ram_reg_116__5_ ( .D(n6298), .CLK(clk), .Q(ram[1861]) );
  DFFPOSX1 ram_reg_116__4_ ( .D(n6297), .CLK(clk), .Q(ram[1860]) );
  DFFPOSX1 ram_reg_116__3_ ( .D(n6296), .CLK(clk), .Q(ram[1859]) );
  DFFPOSX1 ram_reg_116__2_ ( .D(n6295), .CLK(clk), .Q(ram[1858]) );
  DFFPOSX1 ram_reg_116__1_ ( .D(n6294), .CLK(clk), .Q(ram[1857]) );
  DFFPOSX1 ram_reg_116__0_ ( .D(n6293), .CLK(clk), .Q(ram[1856]) );
  DFFPOSX1 ram_reg_115__15_ ( .D(n6292), .CLK(clk), .Q(ram[1855]) );
  DFFPOSX1 ram_reg_115__14_ ( .D(n6291), .CLK(clk), .Q(ram[1854]) );
  DFFPOSX1 ram_reg_115__13_ ( .D(n6290), .CLK(clk), .Q(ram[1853]) );
  DFFPOSX1 ram_reg_115__12_ ( .D(n6289), .CLK(clk), .Q(ram[1852]) );
  DFFPOSX1 ram_reg_115__11_ ( .D(n6288), .CLK(clk), .Q(ram[1851]) );
  DFFPOSX1 ram_reg_115__10_ ( .D(n6287), .CLK(clk), .Q(ram[1850]) );
  DFFPOSX1 ram_reg_115__9_ ( .D(n6286), .CLK(clk), .Q(ram[1849]) );
  DFFPOSX1 ram_reg_115__8_ ( .D(n6285), .CLK(clk), .Q(ram[1848]) );
  DFFPOSX1 ram_reg_115__7_ ( .D(n6284), .CLK(clk), .Q(ram[1847]) );
  DFFPOSX1 ram_reg_115__6_ ( .D(n6283), .CLK(clk), .Q(ram[1846]) );
  DFFPOSX1 ram_reg_115__5_ ( .D(n6282), .CLK(clk), .Q(ram[1845]) );
  DFFPOSX1 ram_reg_115__4_ ( .D(n6281), .CLK(clk), .Q(ram[1844]) );
  DFFPOSX1 ram_reg_115__3_ ( .D(n6280), .CLK(clk), .Q(ram[1843]) );
  DFFPOSX1 ram_reg_115__2_ ( .D(n6279), .CLK(clk), .Q(ram[1842]) );
  DFFPOSX1 ram_reg_115__1_ ( .D(n6278), .CLK(clk), .Q(ram[1841]) );
  DFFPOSX1 ram_reg_115__0_ ( .D(n6277), .CLK(clk), .Q(ram[1840]) );
  DFFPOSX1 ram_reg_114__15_ ( .D(n6276), .CLK(clk), .Q(ram[1839]) );
  DFFPOSX1 ram_reg_114__14_ ( .D(n6275), .CLK(clk), .Q(ram[1838]) );
  DFFPOSX1 ram_reg_114__13_ ( .D(n6274), .CLK(clk), .Q(ram[1837]) );
  DFFPOSX1 ram_reg_114__12_ ( .D(n6273), .CLK(clk), .Q(ram[1836]) );
  DFFPOSX1 ram_reg_114__11_ ( .D(n6272), .CLK(clk), .Q(ram[1835]) );
  DFFPOSX1 ram_reg_114__10_ ( .D(n6271), .CLK(clk), .Q(ram[1834]) );
  DFFPOSX1 ram_reg_114__9_ ( .D(n6270), .CLK(clk), .Q(ram[1833]) );
  DFFPOSX1 ram_reg_114__8_ ( .D(n6269), .CLK(clk), .Q(ram[1832]) );
  DFFPOSX1 ram_reg_114__7_ ( .D(n6268), .CLK(clk), .Q(ram[1831]) );
  DFFPOSX1 ram_reg_114__6_ ( .D(n6267), .CLK(clk), .Q(ram[1830]) );
  DFFPOSX1 ram_reg_114__5_ ( .D(n6266), .CLK(clk), .Q(ram[1829]) );
  DFFPOSX1 ram_reg_114__4_ ( .D(n6265), .CLK(clk), .Q(ram[1828]) );
  DFFPOSX1 ram_reg_114__3_ ( .D(n6264), .CLK(clk), .Q(ram[1827]) );
  DFFPOSX1 ram_reg_114__2_ ( .D(n6263), .CLK(clk), .Q(ram[1826]) );
  DFFPOSX1 ram_reg_114__1_ ( .D(n6262), .CLK(clk), .Q(ram[1825]) );
  DFFPOSX1 ram_reg_114__0_ ( .D(n6261), .CLK(clk), .Q(ram[1824]) );
  DFFPOSX1 ram_reg_113__15_ ( .D(n6260), .CLK(clk), .Q(ram[1823]) );
  DFFPOSX1 ram_reg_113__14_ ( .D(n6259), .CLK(clk), .Q(ram[1822]) );
  DFFPOSX1 ram_reg_113__13_ ( .D(n6258), .CLK(clk), .Q(ram[1821]) );
  DFFPOSX1 ram_reg_113__12_ ( .D(n6257), .CLK(clk), .Q(ram[1820]) );
  DFFPOSX1 ram_reg_113__11_ ( .D(n6256), .CLK(clk), .Q(ram[1819]) );
  DFFPOSX1 ram_reg_113__10_ ( .D(n6255), .CLK(clk), .Q(ram[1818]) );
  DFFPOSX1 ram_reg_113__9_ ( .D(n6254), .CLK(clk), .Q(ram[1817]) );
  DFFPOSX1 ram_reg_113__8_ ( .D(n6253), .CLK(clk), .Q(ram[1816]) );
  DFFPOSX1 ram_reg_113__7_ ( .D(n6252), .CLK(clk), .Q(ram[1815]) );
  DFFPOSX1 ram_reg_113__6_ ( .D(n6251), .CLK(clk), .Q(ram[1814]) );
  DFFPOSX1 ram_reg_113__5_ ( .D(n6250), .CLK(clk), .Q(ram[1813]) );
  DFFPOSX1 ram_reg_113__4_ ( .D(n6249), .CLK(clk), .Q(ram[1812]) );
  DFFPOSX1 ram_reg_113__3_ ( .D(n6248), .CLK(clk), .Q(ram[1811]) );
  DFFPOSX1 ram_reg_113__2_ ( .D(n6247), .CLK(clk), .Q(ram[1810]) );
  DFFPOSX1 ram_reg_113__1_ ( .D(n6246), .CLK(clk), .Q(ram[1809]) );
  DFFPOSX1 ram_reg_113__0_ ( .D(n6245), .CLK(clk), .Q(ram[1808]) );
  DFFPOSX1 ram_reg_112__15_ ( .D(n6244), .CLK(clk), .Q(ram[1807]) );
  DFFPOSX1 ram_reg_112__14_ ( .D(n6243), .CLK(clk), .Q(ram[1806]) );
  DFFPOSX1 ram_reg_112__13_ ( .D(n6242), .CLK(clk), .Q(ram[1805]) );
  DFFPOSX1 ram_reg_112__12_ ( .D(n6241), .CLK(clk), .Q(ram[1804]) );
  DFFPOSX1 ram_reg_112__11_ ( .D(n6240), .CLK(clk), .Q(ram[1803]) );
  DFFPOSX1 ram_reg_112__10_ ( .D(n6239), .CLK(clk), .Q(ram[1802]) );
  DFFPOSX1 ram_reg_112__9_ ( .D(n6238), .CLK(clk), .Q(ram[1801]) );
  DFFPOSX1 ram_reg_112__8_ ( .D(n6237), .CLK(clk), .Q(ram[1800]) );
  DFFPOSX1 ram_reg_112__7_ ( .D(n6236), .CLK(clk), .Q(ram[1799]) );
  DFFPOSX1 ram_reg_112__6_ ( .D(n6235), .CLK(clk), .Q(ram[1798]) );
  DFFPOSX1 ram_reg_112__5_ ( .D(n6234), .CLK(clk), .Q(ram[1797]) );
  DFFPOSX1 ram_reg_112__4_ ( .D(n6233), .CLK(clk), .Q(ram[1796]) );
  DFFPOSX1 ram_reg_112__3_ ( .D(n6232), .CLK(clk), .Q(ram[1795]) );
  DFFPOSX1 ram_reg_112__2_ ( .D(n6231), .CLK(clk), .Q(ram[1794]) );
  DFFPOSX1 ram_reg_112__1_ ( .D(n6230), .CLK(clk), .Q(ram[1793]) );
  DFFPOSX1 ram_reg_112__0_ ( .D(n6229), .CLK(clk), .Q(ram[1792]) );
  DFFPOSX1 ram_reg_111__15_ ( .D(n6228), .CLK(clk), .Q(ram[1791]) );
  DFFPOSX1 ram_reg_111__14_ ( .D(n6227), .CLK(clk), .Q(ram[1790]) );
  DFFPOSX1 ram_reg_111__13_ ( .D(n6226), .CLK(clk), .Q(ram[1789]) );
  DFFPOSX1 ram_reg_111__12_ ( .D(n6225), .CLK(clk), .Q(ram[1788]) );
  DFFPOSX1 ram_reg_111__11_ ( .D(n6224), .CLK(clk), .Q(ram[1787]) );
  DFFPOSX1 ram_reg_111__10_ ( .D(n6223), .CLK(clk), .Q(ram[1786]) );
  DFFPOSX1 ram_reg_111__9_ ( .D(n6222), .CLK(clk), .Q(ram[1785]) );
  DFFPOSX1 ram_reg_111__8_ ( .D(n6221), .CLK(clk), .Q(ram[1784]) );
  DFFPOSX1 ram_reg_111__7_ ( .D(n6220), .CLK(clk), .Q(ram[1783]) );
  DFFPOSX1 ram_reg_111__6_ ( .D(n6219), .CLK(clk), .Q(ram[1782]) );
  DFFPOSX1 ram_reg_111__5_ ( .D(n6218), .CLK(clk), .Q(ram[1781]) );
  DFFPOSX1 ram_reg_111__4_ ( .D(n6217), .CLK(clk), .Q(ram[1780]) );
  DFFPOSX1 ram_reg_111__3_ ( .D(n6216), .CLK(clk), .Q(ram[1779]) );
  DFFPOSX1 ram_reg_111__2_ ( .D(n6215), .CLK(clk), .Q(ram[1778]) );
  DFFPOSX1 ram_reg_111__1_ ( .D(n6214), .CLK(clk), .Q(ram[1777]) );
  DFFPOSX1 ram_reg_111__0_ ( .D(n6213), .CLK(clk), .Q(ram[1776]) );
  DFFPOSX1 ram_reg_110__15_ ( .D(n6212), .CLK(clk), .Q(ram[1775]) );
  DFFPOSX1 ram_reg_110__14_ ( .D(n6211), .CLK(clk), .Q(ram[1774]) );
  DFFPOSX1 ram_reg_110__13_ ( .D(n6210), .CLK(clk), .Q(ram[1773]) );
  DFFPOSX1 ram_reg_110__12_ ( .D(n6209), .CLK(clk), .Q(ram[1772]) );
  DFFPOSX1 ram_reg_110__11_ ( .D(n6208), .CLK(clk), .Q(ram[1771]) );
  DFFPOSX1 ram_reg_110__10_ ( .D(n6207), .CLK(clk), .Q(ram[1770]) );
  DFFPOSX1 ram_reg_110__9_ ( .D(n6206), .CLK(clk), .Q(ram[1769]) );
  DFFPOSX1 ram_reg_110__8_ ( .D(n6205), .CLK(clk), .Q(ram[1768]) );
  DFFPOSX1 ram_reg_110__7_ ( .D(n6204), .CLK(clk), .Q(ram[1767]) );
  DFFPOSX1 ram_reg_110__6_ ( .D(n6203), .CLK(clk), .Q(ram[1766]) );
  DFFPOSX1 ram_reg_110__5_ ( .D(n6202), .CLK(clk), .Q(ram[1765]) );
  DFFPOSX1 ram_reg_110__4_ ( .D(n6201), .CLK(clk), .Q(ram[1764]) );
  DFFPOSX1 ram_reg_110__3_ ( .D(n6200), .CLK(clk), .Q(ram[1763]) );
  DFFPOSX1 ram_reg_110__2_ ( .D(n6199), .CLK(clk), .Q(ram[1762]) );
  DFFPOSX1 ram_reg_110__1_ ( .D(n6198), .CLK(clk), .Q(ram[1761]) );
  DFFPOSX1 ram_reg_110__0_ ( .D(n6197), .CLK(clk), .Q(ram[1760]) );
  DFFPOSX1 ram_reg_109__15_ ( .D(n6196), .CLK(clk), .Q(ram[1759]) );
  DFFPOSX1 ram_reg_109__14_ ( .D(n6195), .CLK(clk), .Q(ram[1758]) );
  DFFPOSX1 ram_reg_109__13_ ( .D(n6194), .CLK(clk), .Q(ram[1757]) );
  DFFPOSX1 ram_reg_109__12_ ( .D(n6193), .CLK(clk), .Q(ram[1756]) );
  DFFPOSX1 ram_reg_109__11_ ( .D(n6192), .CLK(clk), .Q(ram[1755]) );
  DFFPOSX1 ram_reg_109__10_ ( .D(n6191), .CLK(clk), .Q(ram[1754]) );
  DFFPOSX1 ram_reg_109__9_ ( .D(n6190), .CLK(clk), .Q(ram[1753]) );
  DFFPOSX1 ram_reg_109__8_ ( .D(n6189), .CLK(clk), .Q(ram[1752]) );
  DFFPOSX1 ram_reg_109__7_ ( .D(n6188), .CLK(clk), .Q(ram[1751]) );
  DFFPOSX1 ram_reg_109__6_ ( .D(n6187), .CLK(clk), .Q(ram[1750]) );
  DFFPOSX1 ram_reg_109__5_ ( .D(n6186), .CLK(clk), .Q(ram[1749]) );
  DFFPOSX1 ram_reg_109__4_ ( .D(n6185), .CLK(clk), .Q(ram[1748]) );
  DFFPOSX1 ram_reg_109__3_ ( .D(n6184), .CLK(clk), .Q(ram[1747]) );
  DFFPOSX1 ram_reg_109__2_ ( .D(n6183), .CLK(clk), .Q(ram[1746]) );
  DFFPOSX1 ram_reg_109__1_ ( .D(n6182), .CLK(clk), .Q(ram[1745]) );
  DFFPOSX1 ram_reg_109__0_ ( .D(n6181), .CLK(clk), .Q(ram[1744]) );
  DFFPOSX1 ram_reg_108__15_ ( .D(n6180), .CLK(clk), .Q(ram[1743]) );
  DFFPOSX1 ram_reg_108__14_ ( .D(n6179), .CLK(clk), .Q(ram[1742]) );
  DFFPOSX1 ram_reg_108__13_ ( .D(n6178), .CLK(clk), .Q(ram[1741]) );
  DFFPOSX1 ram_reg_108__12_ ( .D(n6177), .CLK(clk), .Q(ram[1740]) );
  DFFPOSX1 ram_reg_108__11_ ( .D(n6176), .CLK(clk), .Q(ram[1739]) );
  DFFPOSX1 ram_reg_108__10_ ( .D(n6175), .CLK(clk), .Q(ram[1738]) );
  DFFPOSX1 ram_reg_108__9_ ( .D(n6174), .CLK(clk), .Q(ram[1737]) );
  DFFPOSX1 ram_reg_108__8_ ( .D(n6173), .CLK(clk), .Q(ram[1736]) );
  DFFPOSX1 ram_reg_108__7_ ( .D(n6172), .CLK(clk), .Q(ram[1735]) );
  DFFPOSX1 ram_reg_108__6_ ( .D(n6171), .CLK(clk), .Q(ram[1734]) );
  DFFPOSX1 ram_reg_108__5_ ( .D(n6170), .CLK(clk), .Q(ram[1733]) );
  DFFPOSX1 ram_reg_108__4_ ( .D(n6169), .CLK(clk), .Q(ram[1732]) );
  DFFPOSX1 ram_reg_108__3_ ( .D(n6168), .CLK(clk), .Q(ram[1731]) );
  DFFPOSX1 ram_reg_108__2_ ( .D(n6167), .CLK(clk), .Q(ram[1730]) );
  DFFPOSX1 ram_reg_108__1_ ( .D(n6166), .CLK(clk), .Q(ram[1729]) );
  DFFPOSX1 ram_reg_108__0_ ( .D(n6165), .CLK(clk), .Q(ram[1728]) );
  DFFPOSX1 ram_reg_107__15_ ( .D(n6164), .CLK(clk), .Q(ram[1727]) );
  DFFPOSX1 ram_reg_107__14_ ( .D(n6163), .CLK(clk), .Q(ram[1726]) );
  DFFPOSX1 ram_reg_107__13_ ( .D(n6162), .CLK(clk), .Q(ram[1725]) );
  DFFPOSX1 ram_reg_107__12_ ( .D(n6161), .CLK(clk), .Q(ram[1724]) );
  DFFPOSX1 ram_reg_107__11_ ( .D(n6160), .CLK(clk), .Q(ram[1723]) );
  DFFPOSX1 ram_reg_107__10_ ( .D(n6159), .CLK(clk), .Q(ram[1722]) );
  DFFPOSX1 ram_reg_107__9_ ( .D(n6158), .CLK(clk), .Q(ram[1721]) );
  DFFPOSX1 ram_reg_107__8_ ( .D(n6157), .CLK(clk), .Q(ram[1720]) );
  DFFPOSX1 ram_reg_107__7_ ( .D(n6156), .CLK(clk), .Q(ram[1719]) );
  DFFPOSX1 ram_reg_107__6_ ( .D(n6155), .CLK(clk), .Q(ram[1718]) );
  DFFPOSX1 ram_reg_107__5_ ( .D(n6154), .CLK(clk), .Q(ram[1717]) );
  DFFPOSX1 ram_reg_107__4_ ( .D(n6153), .CLK(clk), .Q(ram[1716]) );
  DFFPOSX1 ram_reg_107__3_ ( .D(n6152), .CLK(clk), .Q(ram[1715]) );
  DFFPOSX1 ram_reg_107__2_ ( .D(n6151), .CLK(clk), .Q(ram[1714]) );
  DFFPOSX1 ram_reg_107__1_ ( .D(n6150), .CLK(clk), .Q(ram[1713]) );
  DFFPOSX1 ram_reg_107__0_ ( .D(n6149), .CLK(clk), .Q(ram[1712]) );
  DFFPOSX1 ram_reg_106__15_ ( .D(n6148), .CLK(clk), .Q(ram[1711]) );
  DFFPOSX1 ram_reg_106__14_ ( .D(n6147), .CLK(clk), .Q(ram[1710]) );
  DFFPOSX1 ram_reg_106__13_ ( .D(n6146), .CLK(clk), .Q(ram[1709]) );
  DFFPOSX1 ram_reg_106__12_ ( .D(n6145), .CLK(clk), .Q(ram[1708]) );
  DFFPOSX1 ram_reg_106__11_ ( .D(n6144), .CLK(clk), .Q(ram[1707]) );
  DFFPOSX1 ram_reg_106__10_ ( .D(n6143), .CLK(clk), .Q(ram[1706]) );
  DFFPOSX1 ram_reg_106__9_ ( .D(n6142), .CLK(clk), .Q(ram[1705]) );
  DFFPOSX1 ram_reg_106__8_ ( .D(n6141), .CLK(clk), .Q(ram[1704]) );
  DFFPOSX1 ram_reg_106__7_ ( .D(n6140), .CLK(clk), .Q(ram[1703]) );
  DFFPOSX1 ram_reg_106__6_ ( .D(n6139), .CLK(clk), .Q(ram[1702]) );
  DFFPOSX1 ram_reg_106__5_ ( .D(n6138), .CLK(clk), .Q(ram[1701]) );
  DFFPOSX1 ram_reg_106__4_ ( .D(n6137), .CLK(clk), .Q(ram[1700]) );
  DFFPOSX1 ram_reg_106__3_ ( .D(n6136), .CLK(clk), .Q(ram[1699]) );
  DFFPOSX1 ram_reg_106__2_ ( .D(n6135), .CLK(clk), .Q(ram[1698]) );
  DFFPOSX1 ram_reg_106__1_ ( .D(n6134), .CLK(clk), .Q(ram[1697]) );
  DFFPOSX1 ram_reg_106__0_ ( .D(n6133), .CLK(clk), .Q(ram[1696]) );
  DFFPOSX1 ram_reg_105__15_ ( .D(n6132), .CLK(clk), .Q(ram[1695]) );
  DFFPOSX1 ram_reg_105__14_ ( .D(n6131), .CLK(clk), .Q(ram[1694]) );
  DFFPOSX1 ram_reg_105__13_ ( .D(n6130), .CLK(clk), .Q(ram[1693]) );
  DFFPOSX1 ram_reg_105__12_ ( .D(n6129), .CLK(clk), .Q(ram[1692]) );
  DFFPOSX1 ram_reg_105__11_ ( .D(n6128), .CLK(clk), .Q(ram[1691]) );
  DFFPOSX1 ram_reg_105__10_ ( .D(n6127), .CLK(clk), .Q(ram[1690]) );
  DFFPOSX1 ram_reg_105__9_ ( .D(n6126), .CLK(clk), .Q(ram[1689]) );
  DFFPOSX1 ram_reg_105__8_ ( .D(n6125), .CLK(clk), .Q(ram[1688]) );
  DFFPOSX1 ram_reg_105__7_ ( .D(n6124), .CLK(clk), .Q(ram[1687]) );
  DFFPOSX1 ram_reg_105__6_ ( .D(n6123), .CLK(clk), .Q(ram[1686]) );
  DFFPOSX1 ram_reg_105__5_ ( .D(n6122), .CLK(clk), .Q(ram[1685]) );
  DFFPOSX1 ram_reg_105__4_ ( .D(n6121), .CLK(clk), .Q(ram[1684]) );
  DFFPOSX1 ram_reg_105__3_ ( .D(n6120), .CLK(clk), .Q(ram[1683]) );
  DFFPOSX1 ram_reg_105__2_ ( .D(n6119), .CLK(clk), .Q(ram[1682]) );
  DFFPOSX1 ram_reg_105__1_ ( .D(n6118), .CLK(clk), .Q(ram[1681]) );
  DFFPOSX1 ram_reg_105__0_ ( .D(n6117), .CLK(clk), .Q(ram[1680]) );
  DFFPOSX1 ram_reg_104__15_ ( .D(n6116), .CLK(clk), .Q(ram[1679]) );
  DFFPOSX1 ram_reg_104__14_ ( .D(n6115), .CLK(clk), .Q(ram[1678]) );
  DFFPOSX1 ram_reg_104__13_ ( .D(n6114), .CLK(clk), .Q(ram[1677]) );
  DFFPOSX1 ram_reg_104__12_ ( .D(n6113), .CLK(clk), .Q(ram[1676]) );
  DFFPOSX1 ram_reg_104__11_ ( .D(n6112), .CLK(clk), .Q(ram[1675]) );
  DFFPOSX1 ram_reg_104__10_ ( .D(n6111), .CLK(clk), .Q(ram[1674]) );
  DFFPOSX1 ram_reg_104__9_ ( .D(n6110), .CLK(clk), .Q(ram[1673]) );
  DFFPOSX1 ram_reg_104__8_ ( .D(n6109), .CLK(clk), .Q(ram[1672]) );
  DFFPOSX1 ram_reg_104__7_ ( .D(n6108), .CLK(clk), .Q(ram[1671]) );
  DFFPOSX1 ram_reg_104__6_ ( .D(n6107), .CLK(clk), .Q(ram[1670]) );
  DFFPOSX1 ram_reg_104__5_ ( .D(n6106), .CLK(clk), .Q(ram[1669]) );
  DFFPOSX1 ram_reg_104__4_ ( .D(n6105), .CLK(clk), .Q(ram[1668]) );
  DFFPOSX1 ram_reg_104__3_ ( .D(n6104), .CLK(clk), .Q(ram[1667]) );
  DFFPOSX1 ram_reg_104__2_ ( .D(n6103), .CLK(clk), .Q(ram[1666]) );
  DFFPOSX1 ram_reg_104__1_ ( .D(n6102), .CLK(clk), .Q(ram[1665]) );
  DFFPOSX1 ram_reg_104__0_ ( .D(n6101), .CLK(clk), .Q(ram[1664]) );
  DFFPOSX1 ram_reg_103__15_ ( .D(n6100), .CLK(clk), .Q(ram[1663]) );
  DFFPOSX1 ram_reg_103__14_ ( .D(n6099), .CLK(clk), .Q(ram[1662]) );
  DFFPOSX1 ram_reg_103__13_ ( .D(n6098), .CLK(clk), .Q(ram[1661]) );
  DFFPOSX1 ram_reg_103__12_ ( .D(n6097), .CLK(clk), .Q(ram[1660]) );
  DFFPOSX1 ram_reg_103__11_ ( .D(n6096), .CLK(clk), .Q(ram[1659]) );
  DFFPOSX1 ram_reg_103__10_ ( .D(n6095), .CLK(clk), .Q(ram[1658]) );
  DFFPOSX1 ram_reg_103__9_ ( .D(n6094), .CLK(clk), .Q(ram[1657]) );
  DFFPOSX1 ram_reg_103__8_ ( .D(n6093), .CLK(clk), .Q(ram[1656]) );
  DFFPOSX1 ram_reg_103__7_ ( .D(n6092), .CLK(clk), .Q(ram[1655]) );
  DFFPOSX1 ram_reg_103__6_ ( .D(n6091), .CLK(clk), .Q(ram[1654]) );
  DFFPOSX1 ram_reg_103__5_ ( .D(n6090), .CLK(clk), .Q(ram[1653]) );
  DFFPOSX1 ram_reg_103__4_ ( .D(n6089), .CLK(clk), .Q(ram[1652]) );
  DFFPOSX1 ram_reg_103__3_ ( .D(n6088), .CLK(clk), .Q(ram[1651]) );
  DFFPOSX1 ram_reg_103__2_ ( .D(n6087), .CLK(clk), .Q(ram[1650]) );
  DFFPOSX1 ram_reg_103__1_ ( .D(n6086), .CLK(clk), .Q(ram[1649]) );
  DFFPOSX1 ram_reg_103__0_ ( .D(n6085), .CLK(clk), .Q(ram[1648]) );
  DFFPOSX1 ram_reg_102__15_ ( .D(n6084), .CLK(clk), .Q(ram[1647]) );
  DFFPOSX1 ram_reg_102__14_ ( .D(n6083), .CLK(clk), .Q(ram[1646]) );
  DFFPOSX1 ram_reg_102__13_ ( .D(n6082), .CLK(clk), .Q(ram[1645]) );
  DFFPOSX1 ram_reg_102__12_ ( .D(n6081), .CLK(clk), .Q(ram[1644]) );
  DFFPOSX1 ram_reg_102__11_ ( .D(n6080), .CLK(clk), .Q(ram[1643]) );
  DFFPOSX1 ram_reg_102__10_ ( .D(n6079), .CLK(clk), .Q(ram[1642]) );
  DFFPOSX1 ram_reg_102__9_ ( .D(n6078), .CLK(clk), .Q(ram[1641]) );
  DFFPOSX1 ram_reg_102__8_ ( .D(n6077), .CLK(clk), .Q(ram[1640]) );
  DFFPOSX1 ram_reg_102__7_ ( .D(n6076), .CLK(clk), .Q(ram[1639]) );
  DFFPOSX1 ram_reg_102__6_ ( .D(n6075), .CLK(clk), .Q(ram[1638]) );
  DFFPOSX1 ram_reg_102__5_ ( .D(n6074), .CLK(clk), .Q(ram[1637]) );
  DFFPOSX1 ram_reg_102__4_ ( .D(n6073), .CLK(clk), .Q(ram[1636]) );
  DFFPOSX1 ram_reg_102__3_ ( .D(n6072), .CLK(clk), .Q(ram[1635]) );
  DFFPOSX1 ram_reg_102__2_ ( .D(n6071), .CLK(clk), .Q(ram[1634]) );
  DFFPOSX1 ram_reg_102__1_ ( .D(n6070), .CLK(clk), .Q(ram[1633]) );
  DFFPOSX1 ram_reg_102__0_ ( .D(n6069), .CLK(clk), .Q(ram[1632]) );
  DFFPOSX1 ram_reg_101__15_ ( .D(n6068), .CLK(clk), .Q(ram[1631]) );
  DFFPOSX1 ram_reg_101__14_ ( .D(n6067), .CLK(clk), .Q(ram[1630]) );
  DFFPOSX1 ram_reg_101__13_ ( .D(n6066), .CLK(clk), .Q(ram[1629]) );
  DFFPOSX1 ram_reg_101__12_ ( .D(n6065), .CLK(clk), .Q(ram[1628]) );
  DFFPOSX1 ram_reg_101__11_ ( .D(n6064), .CLK(clk), .Q(ram[1627]) );
  DFFPOSX1 ram_reg_101__10_ ( .D(n6063), .CLK(clk), .Q(ram[1626]) );
  DFFPOSX1 ram_reg_101__9_ ( .D(n6062), .CLK(clk), .Q(ram[1625]) );
  DFFPOSX1 ram_reg_101__8_ ( .D(n6061), .CLK(clk), .Q(ram[1624]) );
  DFFPOSX1 ram_reg_101__7_ ( .D(n6060), .CLK(clk), .Q(ram[1623]) );
  DFFPOSX1 ram_reg_101__6_ ( .D(n6059), .CLK(clk), .Q(ram[1622]) );
  DFFPOSX1 ram_reg_101__5_ ( .D(n6058), .CLK(clk), .Q(ram[1621]) );
  DFFPOSX1 ram_reg_101__4_ ( .D(n6057), .CLK(clk), .Q(ram[1620]) );
  DFFPOSX1 ram_reg_101__3_ ( .D(n6056), .CLK(clk), .Q(ram[1619]) );
  DFFPOSX1 ram_reg_101__2_ ( .D(n6055), .CLK(clk), .Q(ram[1618]) );
  DFFPOSX1 ram_reg_101__1_ ( .D(n6054), .CLK(clk), .Q(ram[1617]) );
  DFFPOSX1 ram_reg_101__0_ ( .D(n6053), .CLK(clk), .Q(ram[1616]) );
  DFFPOSX1 ram_reg_100__15_ ( .D(n6052), .CLK(clk), .Q(ram[1615]) );
  DFFPOSX1 ram_reg_100__14_ ( .D(n6051), .CLK(clk), .Q(ram[1614]) );
  DFFPOSX1 ram_reg_100__13_ ( .D(n6050), .CLK(clk), .Q(ram[1613]) );
  DFFPOSX1 ram_reg_100__12_ ( .D(n6049), .CLK(clk), .Q(ram[1612]) );
  DFFPOSX1 ram_reg_100__11_ ( .D(n6048), .CLK(clk), .Q(ram[1611]) );
  DFFPOSX1 ram_reg_100__10_ ( .D(n6047), .CLK(clk), .Q(ram[1610]) );
  DFFPOSX1 ram_reg_100__9_ ( .D(n6046), .CLK(clk), .Q(ram[1609]) );
  DFFPOSX1 ram_reg_100__8_ ( .D(n6045), .CLK(clk), .Q(ram[1608]) );
  DFFPOSX1 ram_reg_100__7_ ( .D(n6044), .CLK(clk), .Q(ram[1607]) );
  DFFPOSX1 ram_reg_100__6_ ( .D(n6043), .CLK(clk), .Q(ram[1606]) );
  DFFPOSX1 ram_reg_100__5_ ( .D(n6042), .CLK(clk), .Q(ram[1605]) );
  DFFPOSX1 ram_reg_100__4_ ( .D(n6041), .CLK(clk), .Q(ram[1604]) );
  DFFPOSX1 ram_reg_100__3_ ( .D(n6040), .CLK(clk), .Q(ram[1603]) );
  DFFPOSX1 ram_reg_100__2_ ( .D(n6039), .CLK(clk), .Q(ram[1602]) );
  DFFPOSX1 ram_reg_100__1_ ( .D(n6038), .CLK(clk), .Q(ram[1601]) );
  DFFPOSX1 ram_reg_100__0_ ( .D(n6037), .CLK(clk), .Q(ram[1600]) );
  DFFPOSX1 ram_reg_99__15_ ( .D(n6036), .CLK(clk), .Q(ram[1599]) );
  DFFPOSX1 ram_reg_99__14_ ( .D(n6035), .CLK(clk), .Q(ram[1598]) );
  DFFPOSX1 ram_reg_99__13_ ( .D(n6034), .CLK(clk), .Q(ram[1597]) );
  DFFPOSX1 ram_reg_99__12_ ( .D(n6033), .CLK(clk), .Q(ram[1596]) );
  DFFPOSX1 ram_reg_99__11_ ( .D(n6032), .CLK(clk), .Q(ram[1595]) );
  DFFPOSX1 ram_reg_99__10_ ( .D(n6031), .CLK(clk), .Q(ram[1594]) );
  DFFPOSX1 ram_reg_99__9_ ( .D(n6030), .CLK(clk), .Q(ram[1593]) );
  DFFPOSX1 ram_reg_99__8_ ( .D(n6029), .CLK(clk), .Q(ram[1592]) );
  DFFPOSX1 ram_reg_99__7_ ( .D(n6028), .CLK(clk), .Q(ram[1591]) );
  DFFPOSX1 ram_reg_99__6_ ( .D(n6027), .CLK(clk), .Q(ram[1590]) );
  DFFPOSX1 ram_reg_99__5_ ( .D(n6026), .CLK(clk), .Q(ram[1589]) );
  DFFPOSX1 ram_reg_99__4_ ( .D(n6025), .CLK(clk), .Q(ram[1588]) );
  DFFPOSX1 ram_reg_99__3_ ( .D(n6024), .CLK(clk), .Q(ram[1587]) );
  DFFPOSX1 ram_reg_99__2_ ( .D(n6023), .CLK(clk), .Q(ram[1586]) );
  DFFPOSX1 ram_reg_99__1_ ( .D(n6022), .CLK(clk), .Q(ram[1585]) );
  DFFPOSX1 ram_reg_99__0_ ( .D(n6021), .CLK(clk), .Q(ram[1584]) );
  DFFPOSX1 ram_reg_98__15_ ( .D(n6020), .CLK(clk), .Q(ram[1583]) );
  DFFPOSX1 ram_reg_98__14_ ( .D(n6019), .CLK(clk), .Q(ram[1582]) );
  DFFPOSX1 ram_reg_98__13_ ( .D(n6018), .CLK(clk), .Q(ram[1581]) );
  DFFPOSX1 ram_reg_98__12_ ( .D(n6017), .CLK(clk), .Q(ram[1580]) );
  DFFPOSX1 ram_reg_98__11_ ( .D(n6016), .CLK(clk), .Q(ram[1579]) );
  DFFPOSX1 ram_reg_98__10_ ( .D(n6015), .CLK(clk), .Q(ram[1578]) );
  DFFPOSX1 ram_reg_98__9_ ( .D(n6014), .CLK(clk), .Q(ram[1577]) );
  DFFPOSX1 ram_reg_98__8_ ( .D(n6013), .CLK(clk), .Q(ram[1576]) );
  DFFPOSX1 ram_reg_98__7_ ( .D(n6012), .CLK(clk), .Q(ram[1575]) );
  DFFPOSX1 ram_reg_98__6_ ( .D(n6011), .CLK(clk), .Q(ram[1574]) );
  DFFPOSX1 ram_reg_98__5_ ( .D(n6010), .CLK(clk), .Q(ram[1573]) );
  DFFPOSX1 ram_reg_98__4_ ( .D(n6009), .CLK(clk), .Q(ram[1572]) );
  DFFPOSX1 ram_reg_98__3_ ( .D(n6008), .CLK(clk), .Q(ram[1571]) );
  DFFPOSX1 ram_reg_98__2_ ( .D(n6007), .CLK(clk), .Q(ram[1570]) );
  DFFPOSX1 ram_reg_98__1_ ( .D(n6006), .CLK(clk), .Q(ram[1569]) );
  DFFPOSX1 ram_reg_98__0_ ( .D(n6005), .CLK(clk), .Q(ram[1568]) );
  DFFPOSX1 ram_reg_97__15_ ( .D(n6004), .CLK(clk), .Q(ram[1567]) );
  DFFPOSX1 ram_reg_97__14_ ( .D(n6003), .CLK(clk), .Q(ram[1566]) );
  DFFPOSX1 ram_reg_97__13_ ( .D(n6002), .CLK(clk), .Q(ram[1565]) );
  DFFPOSX1 ram_reg_97__12_ ( .D(n6001), .CLK(clk), .Q(ram[1564]) );
  DFFPOSX1 ram_reg_97__11_ ( .D(n6000), .CLK(clk), .Q(ram[1563]) );
  DFFPOSX1 ram_reg_97__10_ ( .D(n5999), .CLK(clk), .Q(ram[1562]) );
  DFFPOSX1 ram_reg_97__9_ ( .D(n5998), .CLK(clk), .Q(ram[1561]) );
  DFFPOSX1 ram_reg_97__8_ ( .D(n5997), .CLK(clk), .Q(ram[1560]) );
  DFFPOSX1 ram_reg_97__7_ ( .D(n5996), .CLK(clk), .Q(ram[1559]) );
  DFFPOSX1 ram_reg_97__6_ ( .D(n5995), .CLK(clk), .Q(ram[1558]) );
  DFFPOSX1 ram_reg_97__5_ ( .D(n5994), .CLK(clk), .Q(ram[1557]) );
  DFFPOSX1 ram_reg_97__4_ ( .D(n5993), .CLK(clk), .Q(ram[1556]) );
  DFFPOSX1 ram_reg_97__3_ ( .D(n5992), .CLK(clk), .Q(ram[1555]) );
  DFFPOSX1 ram_reg_97__2_ ( .D(n5991), .CLK(clk), .Q(ram[1554]) );
  DFFPOSX1 ram_reg_97__1_ ( .D(n5990), .CLK(clk), .Q(ram[1553]) );
  DFFPOSX1 ram_reg_97__0_ ( .D(n5989), .CLK(clk), .Q(ram[1552]) );
  DFFPOSX1 ram_reg_96__15_ ( .D(n5988), .CLK(clk), .Q(ram[1551]) );
  DFFPOSX1 ram_reg_96__14_ ( .D(n5987), .CLK(clk), .Q(ram[1550]) );
  DFFPOSX1 ram_reg_96__13_ ( .D(n5986), .CLK(clk), .Q(ram[1549]) );
  DFFPOSX1 ram_reg_96__12_ ( .D(n5985), .CLK(clk), .Q(ram[1548]) );
  DFFPOSX1 ram_reg_96__11_ ( .D(n5984), .CLK(clk), .Q(ram[1547]) );
  DFFPOSX1 ram_reg_96__10_ ( .D(n5983), .CLK(clk), .Q(ram[1546]) );
  DFFPOSX1 ram_reg_96__9_ ( .D(n5982), .CLK(clk), .Q(ram[1545]) );
  DFFPOSX1 ram_reg_96__8_ ( .D(n5981), .CLK(clk), .Q(ram[1544]) );
  DFFPOSX1 ram_reg_96__7_ ( .D(n5980), .CLK(clk), .Q(ram[1543]) );
  DFFPOSX1 ram_reg_96__6_ ( .D(n5979), .CLK(clk), .Q(ram[1542]) );
  DFFPOSX1 ram_reg_96__5_ ( .D(n5978), .CLK(clk), .Q(ram[1541]) );
  DFFPOSX1 ram_reg_96__4_ ( .D(n5977), .CLK(clk), .Q(ram[1540]) );
  DFFPOSX1 ram_reg_96__3_ ( .D(n5976), .CLK(clk), .Q(ram[1539]) );
  DFFPOSX1 ram_reg_96__2_ ( .D(n5975), .CLK(clk), .Q(ram[1538]) );
  DFFPOSX1 ram_reg_96__1_ ( .D(n5974), .CLK(clk), .Q(ram[1537]) );
  DFFPOSX1 ram_reg_96__0_ ( .D(n5973), .CLK(clk), .Q(ram[1536]) );
  DFFPOSX1 ram_reg_95__15_ ( .D(n5972), .CLK(clk), .Q(ram[1535]) );
  DFFPOSX1 ram_reg_95__14_ ( .D(n5971), .CLK(clk), .Q(ram[1534]) );
  DFFPOSX1 ram_reg_95__13_ ( .D(n5970), .CLK(clk), .Q(ram[1533]) );
  DFFPOSX1 ram_reg_95__12_ ( .D(n5969), .CLK(clk), .Q(ram[1532]) );
  DFFPOSX1 ram_reg_95__11_ ( .D(n5968), .CLK(clk), .Q(ram[1531]) );
  DFFPOSX1 ram_reg_95__10_ ( .D(n5967), .CLK(clk), .Q(ram[1530]) );
  DFFPOSX1 ram_reg_95__9_ ( .D(n5966), .CLK(clk), .Q(ram[1529]) );
  DFFPOSX1 ram_reg_95__8_ ( .D(n5965), .CLK(clk), .Q(ram[1528]) );
  DFFPOSX1 ram_reg_95__7_ ( .D(n5964), .CLK(clk), .Q(ram[1527]) );
  DFFPOSX1 ram_reg_95__6_ ( .D(n5963), .CLK(clk), .Q(ram[1526]) );
  DFFPOSX1 ram_reg_95__5_ ( .D(n5962), .CLK(clk), .Q(ram[1525]) );
  DFFPOSX1 ram_reg_95__4_ ( .D(n5961), .CLK(clk), .Q(ram[1524]) );
  DFFPOSX1 ram_reg_95__3_ ( .D(n5960), .CLK(clk), .Q(ram[1523]) );
  DFFPOSX1 ram_reg_95__2_ ( .D(n5959), .CLK(clk), .Q(ram[1522]) );
  DFFPOSX1 ram_reg_95__1_ ( .D(n5958), .CLK(clk), .Q(ram[1521]) );
  DFFPOSX1 ram_reg_95__0_ ( .D(n5957), .CLK(clk), .Q(ram[1520]) );
  DFFPOSX1 ram_reg_94__15_ ( .D(n5956), .CLK(clk), .Q(ram[1519]) );
  DFFPOSX1 ram_reg_94__14_ ( .D(n5955), .CLK(clk), .Q(ram[1518]) );
  DFFPOSX1 ram_reg_94__13_ ( .D(n5954), .CLK(clk), .Q(ram[1517]) );
  DFFPOSX1 ram_reg_94__12_ ( .D(n5953), .CLK(clk), .Q(ram[1516]) );
  DFFPOSX1 ram_reg_94__11_ ( .D(n5952), .CLK(clk), .Q(ram[1515]) );
  DFFPOSX1 ram_reg_94__10_ ( .D(n5951), .CLK(clk), .Q(ram[1514]) );
  DFFPOSX1 ram_reg_94__9_ ( .D(n5950), .CLK(clk), .Q(ram[1513]) );
  DFFPOSX1 ram_reg_94__8_ ( .D(n5949), .CLK(clk), .Q(ram[1512]) );
  DFFPOSX1 ram_reg_94__7_ ( .D(n5948), .CLK(clk), .Q(ram[1511]) );
  DFFPOSX1 ram_reg_94__6_ ( .D(n5947), .CLK(clk), .Q(ram[1510]) );
  DFFPOSX1 ram_reg_94__5_ ( .D(n5946), .CLK(clk), .Q(ram[1509]) );
  DFFPOSX1 ram_reg_94__4_ ( .D(n5945), .CLK(clk), .Q(ram[1508]) );
  DFFPOSX1 ram_reg_94__3_ ( .D(n5944), .CLK(clk), .Q(ram[1507]) );
  DFFPOSX1 ram_reg_94__2_ ( .D(n5943), .CLK(clk), .Q(ram[1506]) );
  DFFPOSX1 ram_reg_94__1_ ( .D(n5942), .CLK(clk), .Q(ram[1505]) );
  DFFPOSX1 ram_reg_94__0_ ( .D(n5941), .CLK(clk), .Q(ram[1504]) );
  DFFPOSX1 ram_reg_93__15_ ( .D(n5940), .CLK(clk), .Q(ram[1503]) );
  DFFPOSX1 ram_reg_93__14_ ( .D(n5939), .CLK(clk), .Q(ram[1502]) );
  DFFPOSX1 ram_reg_93__13_ ( .D(n5938), .CLK(clk), .Q(ram[1501]) );
  DFFPOSX1 ram_reg_93__12_ ( .D(n5937), .CLK(clk), .Q(ram[1500]) );
  DFFPOSX1 ram_reg_93__11_ ( .D(n5936), .CLK(clk), .Q(ram[1499]) );
  DFFPOSX1 ram_reg_93__10_ ( .D(n5935), .CLK(clk), .Q(ram[1498]) );
  DFFPOSX1 ram_reg_93__9_ ( .D(n5934), .CLK(clk), .Q(ram[1497]) );
  DFFPOSX1 ram_reg_93__8_ ( .D(n5933), .CLK(clk), .Q(ram[1496]) );
  DFFPOSX1 ram_reg_93__7_ ( .D(n5932), .CLK(clk), .Q(ram[1495]) );
  DFFPOSX1 ram_reg_93__6_ ( .D(n5931), .CLK(clk), .Q(ram[1494]) );
  DFFPOSX1 ram_reg_93__5_ ( .D(n5930), .CLK(clk), .Q(ram[1493]) );
  DFFPOSX1 ram_reg_93__4_ ( .D(n5929), .CLK(clk), .Q(ram[1492]) );
  DFFPOSX1 ram_reg_93__3_ ( .D(n5928), .CLK(clk), .Q(ram[1491]) );
  DFFPOSX1 ram_reg_93__2_ ( .D(n5927), .CLK(clk), .Q(ram[1490]) );
  DFFPOSX1 ram_reg_93__1_ ( .D(n5926), .CLK(clk), .Q(ram[1489]) );
  DFFPOSX1 ram_reg_93__0_ ( .D(n5925), .CLK(clk), .Q(ram[1488]) );
  DFFPOSX1 ram_reg_92__15_ ( .D(n5924), .CLK(clk), .Q(ram[1487]) );
  DFFPOSX1 ram_reg_92__14_ ( .D(n5923), .CLK(clk), .Q(ram[1486]) );
  DFFPOSX1 ram_reg_92__13_ ( .D(n5922), .CLK(clk), .Q(ram[1485]) );
  DFFPOSX1 ram_reg_92__12_ ( .D(n5921), .CLK(clk), .Q(ram[1484]) );
  DFFPOSX1 ram_reg_92__11_ ( .D(n5920), .CLK(clk), .Q(ram[1483]) );
  DFFPOSX1 ram_reg_92__10_ ( .D(n5919), .CLK(clk), .Q(ram[1482]) );
  DFFPOSX1 ram_reg_92__9_ ( .D(n5918), .CLK(clk), .Q(ram[1481]) );
  DFFPOSX1 ram_reg_92__8_ ( .D(n5917), .CLK(clk), .Q(ram[1480]) );
  DFFPOSX1 ram_reg_92__7_ ( .D(n5916), .CLK(clk), .Q(ram[1479]) );
  DFFPOSX1 ram_reg_92__6_ ( .D(n5915), .CLK(clk), .Q(ram[1478]) );
  DFFPOSX1 ram_reg_92__5_ ( .D(n5914), .CLK(clk), .Q(ram[1477]) );
  DFFPOSX1 ram_reg_92__4_ ( .D(n5913), .CLK(clk), .Q(ram[1476]) );
  DFFPOSX1 ram_reg_92__3_ ( .D(n5912), .CLK(clk), .Q(ram[1475]) );
  DFFPOSX1 ram_reg_92__2_ ( .D(n5911), .CLK(clk), .Q(ram[1474]) );
  DFFPOSX1 ram_reg_92__1_ ( .D(n5910), .CLK(clk), .Q(ram[1473]) );
  DFFPOSX1 ram_reg_92__0_ ( .D(n5909), .CLK(clk), .Q(ram[1472]) );
  DFFPOSX1 ram_reg_91__15_ ( .D(n5908), .CLK(clk), .Q(ram[1471]) );
  DFFPOSX1 ram_reg_91__14_ ( .D(n5907), .CLK(clk), .Q(ram[1470]) );
  DFFPOSX1 ram_reg_91__13_ ( .D(n5906), .CLK(clk), .Q(ram[1469]) );
  DFFPOSX1 ram_reg_91__12_ ( .D(n5905), .CLK(clk), .Q(ram[1468]) );
  DFFPOSX1 ram_reg_91__11_ ( .D(n5904), .CLK(clk), .Q(ram[1467]) );
  DFFPOSX1 ram_reg_91__10_ ( .D(n5903), .CLK(clk), .Q(ram[1466]) );
  DFFPOSX1 ram_reg_91__9_ ( .D(n5902), .CLK(clk), .Q(ram[1465]) );
  DFFPOSX1 ram_reg_91__8_ ( .D(n5901), .CLK(clk), .Q(ram[1464]) );
  DFFPOSX1 ram_reg_91__7_ ( .D(n5900), .CLK(clk), .Q(ram[1463]) );
  DFFPOSX1 ram_reg_91__6_ ( .D(n5899), .CLK(clk), .Q(ram[1462]) );
  DFFPOSX1 ram_reg_91__5_ ( .D(n5898), .CLK(clk), .Q(ram[1461]) );
  DFFPOSX1 ram_reg_91__4_ ( .D(n5897), .CLK(clk), .Q(ram[1460]) );
  DFFPOSX1 ram_reg_91__3_ ( .D(n5896), .CLK(clk), .Q(ram[1459]) );
  DFFPOSX1 ram_reg_91__2_ ( .D(n5895), .CLK(clk), .Q(ram[1458]) );
  DFFPOSX1 ram_reg_91__1_ ( .D(n5894), .CLK(clk), .Q(ram[1457]) );
  DFFPOSX1 ram_reg_91__0_ ( .D(n5893), .CLK(clk), .Q(ram[1456]) );
  DFFPOSX1 ram_reg_90__15_ ( .D(n5892), .CLK(clk), .Q(ram[1455]) );
  DFFPOSX1 ram_reg_90__14_ ( .D(n5891), .CLK(clk), .Q(ram[1454]) );
  DFFPOSX1 ram_reg_90__13_ ( .D(n5890), .CLK(clk), .Q(ram[1453]) );
  DFFPOSX1 ram_reg_90__12_ ( .D(n5889), .CLK(clk), .Q(ram[1452]) );
  DFFPOSX1 ram_reg_90__11_ ( .D(n5888), .CLK(clk), .Q(ram[1451]) );
  DFFPOSX1 ram_reg_90__10_ ( .D(n5887), .CLK(clk), .Q(ram[1450]) );
  DFFPOSX1 ram_reg_90__9_ ( .D(n5886), .CLK(clk), .Q(ram[1449]) );
  DFFPOSX1 ram_reg_90__8_ ( .D(n5885), .CLK(clk), .Q(ram[1448]) );
  DFFPOSX1 ram_reg_90__7_ ( .D(n5884), .CLK(clk), .Q(ram[1447]) );
  DFFPOSX1 ram_reg_90__6_ ( .D(n5883), .CLK(clk), .Q(ram[1446]) );
  DFFPOSX1 ram_reg_90__5_ ( .D(n5882), .CLK(clk), .Q(ram[1445]) );
  DFFPOSX1 ram_reg_90__4_ ( .D(n5881), .CLK(clk), .Q(ram[1444]) );
  DFFPOSX1 ram_reg_90__3_ ( .D(n5880), .CLK(clk), .Q(ram[1443]) );
  DFFPOSX1 ram_reg_90__2_ ( .D(n5879), .CLK(clk), .Q(ram[1442]) );
  DFFPOSX1 ram_reg_90__1_ ( .D(n5878), .CLK(clk), .Q(ram[1441]) );
  DFFPOSX1 ram_reg_90__0_ ( .D(n5877), .CLK(clk), .Q(ram[1440]) );
  DFFPOSX1 ram_reg_89__15_ ( .D(n5876), .CLK(clk), .Q(ram[1439]) );
  DFFPOSX1 ram_reg_89__14_ ( .D(n5875), .CLK(clk), .Q(ram[1438]) );
  DFFPOSX1 ram_reg_89__13_ ( .D(n5874), .CLK(clk), .Q(ram[1437]) );
  DFFPOSX1 ram_reg_89__12_ ( .D(n5873), .CLK(clk), .Q(ram[1436]) );
  DFFPOSX1 ram_reg_89__11_ ( .D(n5872), .CLK(clk), .Q(ram[1435]) );
  DFFPOSX1 ram_reg_89__10_ ( .D(n5871), .CLK(clk), .Q(ram[1434]) );
  DFFPOSX1 ram_reg_89__9_ ( .D(n5870), .CLK(clk), .Q(ram[1433]) );
  DFFPOSX1 ram_reg_89__8_ ( .D(n5869), .CLK(clk), .Q(ram[1432]) );
  DFFPOSX1 ram_reg_89__7_ ( .D(n5868), .CLK(clk), .Q(ram[1431]) );
  DFFPOSX1 ram_reg_89__6_ ( .D(n5867), .CLK(clk), .Q(ram[1430]) );
  DFFPOSX1 ram_reg_89__5_ ( .D(n5866), .CLK(clk), .Q(ram[1429]) );
  DFFPOSX1 ram_reg_89__4_ ( .D(n5865), .CLK(clk), .Q(ram[1428]) );
  DFFPOSX1 ram_reg_89__3_ ( .D(n5864), .CLK(clk), .Q(ram[1427]) );
  DFFPOSX1 ram_reg_89__2_ ( .D(n5863), .CLK(clk), .Q(ram[1426]) );
  DFFPOSX1 ram_reg_89__1_ ( .D(n5862), .CLK(clk), .Q(ram[1425]) );
  DFFPOSX1 ram_reg_89__0_ ( .D(n5861), .CLK(clk), .Q(ram[1424]) );
  DFFPOSX1 ram_reg_88__15_ ( .D(n5860), .CLK(clk), .Q(ram[1423]) );
  DFFPOSX1 ram_reg_88__14_ ( .D(n5859), .CLK(clk), .Q(ram[1422]) );
  DFFPOSX1 ram_reg_88__13_ ( .D(n5858), .CLK(clk), .Q(ram[1421]) );
  DFFPOSX1 ram_reg_88__12_ ( .D(n5857), .CLK(clk), .Q(ram[1420]) );
  DFFPOSX1 ram_reg_88__11_ ( .D(n5856), .CLK(clk), .Q(ram[1419]) );
  DFFPOSX1 ram_reg_88__10_ ( .D(n5855), .CLK(clk), .Q(ram[1418]) );
  DFFPOSX1 ram_reg_88__9_ ( .D(n5854), .CLK(clk), .Q(ram[1417]) );
  DFFPOSX1 ram_reg_88__8_ ( .D(n5853), .CLK(clk), .Q(ram[1416]) );
  DFFPOSX1 ram_reg_88__7_ ( .D(n5852), .CLK(clk), .Q(ram[1415]) );
  DFFPOSX1 ram_reg_88__6_ ( .D(n5851), .CLK(clk), .Q(ram[1414]) );
  DFFPOSX1 ram_reg_88__5_ ( .D(n5850), .CLK(clk), .Q(ram[1413]) );
  DFFPOSX1 ram_reg_88__4_ ( .D(n5849), .CLK(clk), .Q(ram[1412]) );
  DFFPOSX1 ram_reg_88__3_ ( .D(n5848), .CLK(clk), .Q(ram[1411]) );
  DFFPOSX1 ram_reg_88__2_ ( .D(n5847), .CLK(clk), .Q(ram[1410]) );
  DFFPOSX1 ram_reg_88__1_ ( .D(n5846), .CLK(clk), .Q(ram[1409]) );
  DFFPOSX1 ram_reg_88__0_ ( .D(n5845), .CLK(clk), .Q(ram[1408]) );
  DFFPOSX1 ram_reg_87__15_ ( .D(n5844), .CLK(clk), .Q(ram[1407]) );
  DFFPOSX1 ram_reg_87__14_ ( .D(n5843), .CLK(clk), .Q(ram[1406]) );
  DFFPOSX1 ram_reg_87__13_ ( .D(n5842), .CLK(clk), .Q(ram[1405]) );
  DFFPOSX1 ram_reg_87__12_ ( .D(n5841), .CLK(clk), .Q(ram[1404]) );
  DFFPOSX1 ram_reg_87__11_ ( .D(n5840), .CLK(clk), .Q(ram[1403]) );
  DFFPOSX1 ram_reg_87__10_ ( .D(n5839), .CLK(clk), .Q(ram[1402]) );
  DFFPOSX1 ram_reg_87__9_ ( .D(n5838), .CLK(clk), .Q(ram[1401]) );
  DFFPOSX1 ram_reg_87__8_ ( .D(n5837), .CLK(clk), .Q(ram[1400]) );
  DFFPOSX1 ram_reg_87__7_ ( .D(n5836), .CLK(clk), .Q(ram[1399]) );
  DFFPOSX1 ram_reg_87__6_ ( .D(n5835), .CLK(clk), .Q(ram[1398]) );
  DFFPOSX1 ram_reg_87__5_ ( .D(n5834), .CLK(clk), .Q(ram[1397]) );
  DFFPOSX1 ram_reg_87__4_ ( .D(n5833), .CLK(clk), .Q(ram[1396]) );
  DFFPOSX1 ram_reg_87__3_ ( .D(n5832), .CLK(clk), .Q(ram[1395]) );
  DFFPOSX1 ram_reg_87__2_ ( .D(n5831), .CLK(clk), .Q(ram[1394]) );
  DFFPOSX1 ram_reg_87__1_ ( .D(n5830), .CLK(clk), .Q(ram[1393]) );
  DFFPOSX1 ram_reg_87__0_ ( .D(n5829), .CLK(clk), .Q(ram[1392]) );
  DFFPOSX1 ram_reg_86__15_ ( .D(n5828), .CLK(clk), .Q(ram[1391]) );
  DFFPOSX1 ram_reg_86__14_ ( .D(n5827), .CLK(clk), .Q(ram[1390]) );
  DFFPOSX1 ram_reg_86__13_ ( .D(n5826), .CLK(clk), .Q(ram[1389]) );
  DFFPOSX1 ram_reg_86__12_ ( .D(n5825), .CLK(clk), .Q(ram[1388]) );
  DFFPOSX1 ram_reg_86__11_ ( .D(n5824), .CLK(clk), .Q(ram[1387]) );
  DFFPOSX1 ram_reg_86__10_ ( .D(n5823), .CLK(clk), .Q(ram[1386]) );
  DFFPOSX1 ram_reg_86__9_ ( .D(n5822), .CLK(clk), .Q(ram[1385]) );
  DFFPOSX1 ram_reg_86__8_ ( .D(n5821), .CLK(clk), .Q(ram[1384]) );
  DFFPOSX1 ram_reg_86__7_ ( .D(n5820), .CLK(clk), .Q(ram[1383]) );
  DFFPOSX1 ram_reg_86__6_ ( .D(n5819), .CLK(clk), .Q(ram[1382]) );
  DFFPOSX1 ram_reg_86__5_ ( .D(n5818), .CLK(clk), .Q(ram[1381]) );
  DFFPOSX1 ram_reg_86__4_ ( .D(n5817), .CLK(clk), .Q(ram[1380]) );
  DFFPOSX1 ram_reg_86__3_ ( .D(n5816), .CLK(clk), .Q(ram[1379]) );
  DFFPOSX1 ram_reg_86__2_ ( .D(n5815), .CLK(clk), .Q(ram[1378]) );
  DFFPOSX1 ram_reg_86__1_ ( .D(n5814), .CLK(clk), .Q(ram[1377]) );
  DFFPOSX1 ram_reg_86__0_ ( .D(n5813), .CLK(clk), .Q(ram[1376]) );
  DFFPOSX1 ram_reg_85__15_ ( .D(n5812), .CLK(clk), .Q(ram[1375]) );
  DFFPOSX1 ram_reg_85__14_ ( .D(n5811), .CLK(clk), .Q(ram[1374]) );
  DFFPOSX1 ram_reg_85__13_ ( .D(n5810), .CLK(clk), .Q(ram[1373]) );
  DFFPOSX1 ram_reg_85__12_ ( .D(n5809), .CLK(clk), .Q(ram[1372]) );
  DFFPOSX1 ram_reg_85__11_ ( .D(n5808), .CLK(clk), .Q(ram[1371]) );
  DFFPOSX1 ram_reg_85__10_ ( .D(n5807), .CLK(clk), .Q(ram[1370]) );
  DFFPOSX1 ram_reg_85__9_ ( .D(n5806), .CLK(clk), .Q(ram[1369]) );
  DFFPOSX1 ram_reg_85__8_ ( .D(n5805), .CLK(clk), .Q(ram[1368]) );
  DFFPOSX1 ram_reg_85__7_ ( .D(n5804), .CLK(clk), .Q(ram[1367]) );
  DFFPOSX1 ram_reg_85__6_ ( .D(n5803), .CLK(clk), .Q(ram[1366]) );
  DFFPOSX1 ram_reg_85__5_ ( .D(n5802), .CLK(clk), .Q(ram[1365]) );
  DFFPOSX1 ram_reg_85__4_ ( .D(n5801), .CLK(clk), .Q(ram[1364]) );
  DFFPOSX1 ram_reg_85__3_ ( .D(n5800), .CLK(clk), .Q(ram[1363]) );
  DFFPOSX1 ram_reg_85__2_ ( .D(n5799), .CLK(clk), .Q(ram[1362]) );
  DFFPOSX1 ram_reg_85__1_ ( .D(n5798), .CLK(clk), .Q(ram[1361]) );
  DFFPOSX1 ram_reg_85__0_ ( .D(n5797), .CLK(clk), .Q(ram[1360]) );
  DFFPOSX1 ram_reg_84__15_ ( .D(n5796), .CLK(clk), .Q(ram[1359]) );
  DFFPOSX1 ram_reg_84__14_ ( .D(n5795), .CLK(clk), .Q(ram[1358]) );
  DFFPOSX1 ram_reg_84__13_ ( .D(n5794), .CLK(clk), .Q(ram[1357]) );
  DFFPOSX1 ram_reg_84__12_ ( .D(n5793), .CLK(clk), .Q(ram[1356]) );
  DFFPOSX1 ram_reg_84__11_ ( .D(n5792), .CLK(clk), .Q(ram[1355]) );
  DFFPOSX1 ram_reg_84__10_ ( .D(n5791), .CLK(clk), .Q(ram[1354]) );
  DFFPOSX1 ram_reg_84__9_ ( .D(n5790), .CLK(clk), .Q(ram[1353]) );
  DFFPOSX1 ram_reg_84__8_ ( .D(n5789), .CLK(clk), .Q(ram[1352]) );
  DFFPOSX1 ram_reg_84__7_ ( .D(n5788), .CLK(clk), .Q(ram[1351]) );
  DFFPOSX1 ram_reg_84__6_ ( .D(n5787), .CLK(clk), .Q(ram[1350]) );
  DFFPOSX1 ram_reg_84__5_ ( .D(n5786), .CLK(clk), .Q(ram[1349]) );
  DFFPOSX1 ram_reg_84__4_ ( .D(n5785), .CLK(clk), .Q(ram[1348]) );
  DFFPOSX1 ram_reg_84__3_ ( .D(n5784), .CLK(clk), .Q(ram[1347]) );
  DFFPOSX1 ram_reg_84__2_ ( .D(n5783), .CLK(clk), .Q(ram[1346]) );
  DFFPOSX1 ram_reg_84__1_ ( .D(n5782), .CLK(clk), .Q(ram[1345]) );
  DFFPOSX1 ram_reg_84__0_ ( .D(n5781), .CLK(clk), .Q(ram[1344]) );
  DFFPOSX1 ram_reg_83__15_ ( .D(n5780), .CLK(clk), .Q(ram[1343]) );
  DFFPOSX1 ram_reg_83__14_ ( .D(n5779), .CLK(clk), .Q(ram[1342]) );
  DFFPOSX1 ram_reg_83__13_ ( .D(n5778), .CLK(clk), .Q(ram[1341]) );
  DFFPOSX1 ram_reg_83__12_ ( .D(n5777), .CLK(clk), .Q(ram[1340]) );
  DFFPOSX1 ram_reg_83__11_ ( .D(n5776), .CLK(clk), .Q(ram[1339]) );
  DFFPOSX1 ram_reg_83__10_ ( .D(n5775), .CLK(clk), .Q(ram[1338]) );
  DFFPOSX1 ram_reg_83__9_ ( .D(n5774), .CLK(clk), .Q(ram[1337]) );
  DFFPOSX1 ram_reg_83__8_ ( .D(n5773), .CLK(clk), .Q(ram[1336]) );
  DFFPOSX1 ram_reg_83__7_ ( .D(n5772), .CLK(clk), .Q(ram[1335]) );
  DFFPOSX1 ram_reg_83__6_ ( .D(n5771), .CLK(clk), .Q(ram[1334]) );
  DFFPOSX1 ram_reg_83__5_ ( .D(n5770), .CLK(clk), .Q(ram[1333]) );
  DFFPOSX1 ram_reg_83__4_ ( .D(n5769), .CLK(clk), .Q(ram[1332]) );
  DFFPOSX1 ram_reg_83__3_ ( .D(n5768), .CLK(clk), .Q(ram[1331]) );
  DFFPOSX1 ram_reg_83__2_ ( .D(n5767), .CLK(clk), .Q(ram[1330]) );
  DFFPOSX1 ram_reg_83__1_ ( .D(n5766), .CLK(clk), .Q(ram[1329]) );
  DFFPOSX1 ram_reg_83__0_ ( .D(n5765), .CLK(clk), .Q(ram[1328]) );
  DFFPOSX1 ram_reg_82__15_ ( .D(n5764), .CLK(clk), .Q(ram[1327]) );
  DFFPOSX1 ram_reg_82__14_ ( .D(n5763), .CLK(clk), .Q(ram[1326]) );
  DFFPOSX1 ram_reg_82__13_ ( .D(n5762), .CLK(clk), .Q(ram[1325]) );
  DFFPOSX1 ram_reg_82__12_ ( .D(n5761), .CLK(clk), .Q(ram[1324]) );
  DFFPOSX1 ram_reg_82__11_ ( .D(n5760), .CLK(clk), .Q(ram[1323]) );
  DFFPOSX1 ram_reg_82__10_ ( .D(n5759), .CLK(clk), .Q(ram[1322]) );
  DFFPOSX1 ram_reg_82__9_ ( .D(n5758), .CLK(clk), .Q(ram[1321]) );
  DFFPOSX1 ram_reg_82__8_ ( .D(n5757), .CLK(clk), .Q(ram[1320]) );
  DFFPOSX1 ram_reg_82__7_ ( .D(n5756), .CLK(clk), .Q(ram[1319]) );
  DFFPOSX1 ram_reg_82__6_ ( .D(n5755), .CLK(clk), .Q(ram[1318]) );
  DFFPOSX1 ram_reg_82__5_ ( .D(n5754), .CLK(clk), .Q(ram[1317]) );
  DFFPOSX1 ram_reg_82__4_ ( .D(n5753), .CLK(clk), .Q(ram[1316]) );
  DFFPOSX1 ram_reg_82__3_ ( .D(n5752), .CLK(clk), .Q(ram[1315]) );
  DFFPOSX1 ram_reg_82__2_ ( .D(n5751), .CLK(clk), .Q(ram[1314]) );
  DFFPOSX1 ram_reg_82__1_ ( .D(n5750), .CLK(clk), .Q(ram[1313]) );
  DFFPOSX1 ram_reg_82__0_ ( .D(n5749), .CLK(clk), .Q(ram[1312]) );
  DFFPOSX1 ram_reg_81__15_ ( .D(n5748), .CLK(clk), .Q(ram[1311]) );
  DFFPOSX1 ram_reg_81__14_ ( .D(n5747), .CLK(clk), .Q(ram[1310]) );
  DFFPOSX1 ram_reg_81__13_ ( .D(n5746), .CLK(clk), .Q(ram[1309]) );
  DFFPOSX1 ram_reg_81__12_ ( .D(n5745), .CLK(clk), .Q(ram[1308]) );
  DFFPOSX1 ram_reg_81__11_ ( .D(n5744), .CLK(clk), .Q(ram[1307]) );
  DFFPOSX1 ram_reg_81__10_ ( .D(n5743), .CLK(clk), .Q(ram[1306]) );
  DFFPOSX1 ram_reg_81__9_ ( .D(n5742), .CLK(clk), .Q(ram[1305]) );
  DFFPOSX1 ram_reg_81__8_ ( .D(n5741), .CLK(clk), .Q(ram[1304]) );
  DFFPOSX1 ram_reg_81__7_ ( .D(n5740), .CLK(clk), .Q(ram[1303]) );
  DFFPOSX1 ram_reg_81__6_ ( .D(n5739), .CLK(clk), .Q(ram[1302]) );
  DFFPOSX1 ram_reg_81__5_ ( .D(n5738), .CLK(clk), .Q(ram[1301]) );
  DFFPOSX1 ram_reg_81__4_ ( .D(n5737), .CLK(clk), .Q(ram[1300]) );
  DFFPOSX1 ram_reg_81__3_ ( .D(n5736), .CLK(clk), .Q(ram[1299]) );
  DFFPOSX1 ram_reg_81__2_ ( .D(n5735), .CLK(clk), .Q(ram[1298]) );
  DFFPOSX1 ram_reg_81__1_ ( .D(n5734), .CLK(clk), .Q(ram[1297]) );
  DFFPOSX1 ram_reg_81__0_ ( .D(n5733), .CLK(clk), .Q(ram[1296]) );
  DFFPOSX1 ram_reg_80__15_ ( .D(n5732), .CLK(clk), .Q(ram[1295]) );
  DFFPOSX1 ram_reg_80__14_ ( .D(n5731), .CLK(clk), .Q(ram[1294]) );
  DFFPOSX1 ram_reg_80__13_ ( .D(n5730), .CLK(clk), .Q(ram[1293]) );
  DFFPOSX1 ram_reg_80__12_ ( .D(n5729), .CLK(clk), .Q(ram[1292]) );
  DFFPOSX1 ram_reg_80__11_ ( .D(n5728), .CLK(clk), .Q(ram[1291]) );
  DFFPOSX1 ram_reg_80__10_ ( .D(n5727), .CLK(clk), .Q(ram[1290]) );
  DFFPOSX1 ram_reg_80__9_ ( .D(n5726), .CLK(clk), .Q(ram[1289]) );
  DFFPOSX1 ram_reg_80__8_ ( .D(n5725), .CLK(clk), .Q(ram[1288]) );
  DFFPOSX1 ram_reg_80__7_ ( .D(n5724), .CLK(clk), .Q(ram[1287]) );
  DFFPOSX1 ram_reg_80__6_ ( .D(n5723), .CLK(clk), .Q(ram[1286]) );
  DFFPOSX1 ram_reg_80__5_ ( .D(n5722), .CLK(clk), .Q(ram[1285]) );
  DFFPOSX1 ram_reg_80__4_ ( .D(n5721), .CLK(clk), .Q(ram[1284]) );
  DFFPOSX1 ram_reg_80__3_ ( .D(n5720), .CLK(clk), .Q(ram[1283]) );
  DFFPOSX1 ram_reg_80__2_ ( .D(n5719), .CLK(clk), .Q(ram[1282]) );
  DFFPOSX1 ram_reg_80__1_ ( .D(n5718), .CLK(clk), .Q(ram[1281]) );
  DFFPOSX1 ram_reg_80__0_ ( .D(n5717), .CLK(clk), .Q(ram[1280]) );
  DFFPOSX1 ram_reg_79__15_ ( .D(n5716), .CLK(clk), .Q(ram[1279]) );
  DFFPOSX1 ram_reg_79__14_ ( .D(n5715), .CLK(clk), .Q(ram[1278]) );
  DFFPOSX1 ram_reg_79__13_ ( .D(n5714), .CLK(clk), .Q(ram[1277]) );
  DFFPOSX1 ram_reg_79__12_ ( .D(n5713), .CLK(clk), .Q(ram[1276]) );
  DFFPOSX1 ram_reg_79__11_ ( .D(n5712), .CLK(clk), .Q(ram[1275]) );
  DFFPOSX1 ram_reg_79__10_ ( .D(n5711), .CLK(clk), .Q(ram[1274]) );
  DFFPOSX1 ram_reg_79__9_ ( .D(n5710), .CLK(clk), .Q(ram[1273]) );
  DFFPOSX1 ram_reg_79__8_ ( .D(n5709), .CLK(clk), .Q(ram[1272]) );
  DFFPOSX1 ram_reg_79__7_ ( .D(n5708), .CLK(clk), .Q(ram[1271]) );
  DFFPOSX1 ram_reg_79__6_ ( .D(n5707), .CLK(clk), .Q(ram[1270]) );
  DFFPOSX1 ram_reg_79__5_ ( .D(n5706), .CLK(clk), .Q(ram[1269]) );
  DFFPOSX1 ram_reg_79__4_ ( .D(n5705), .CLK(clk), .Q(ram[1268]) );
  DFFPOSX1 ram_reg_79__3_ ( .D(n5704), .CLK(clk), .Q(ram[1267]) );
  DFFPOSX1 ram_reg_79__2_ ( .D(n5703), .CLK(clk), .Q(ram[1266]) );
  DFFPOSX1 ram_reg_79__1_ ( .D(n5702), .CLK(clk), .Q(ram[1265]) );
  DFFPOSX1 ram_reg_79__0_ ( .D(n5701), .CLK(clk), .Q(ram[1264]) );
  DFFPOSX1 ram_reg_78__15_ ( .D(n5700), .CLK(clk), .Q(ram[1263]) );
  DFFPOSX1 ram_reg_78__14_ ( .D(n5699), .CLK(clk), .Q(ram[1262]) );
  DFFPOSX1 ram_reg_78__13_ ( .D(n5698), .CLK(clk), .Q(ram[1261]) );
  DFFPOSX1 ram_reg_78__12_ ( .D(n5697), .CLK(clk), .Q(ram[1260]) );
  DFFPOSX1 ram_reg_78__11_ ( .D(n5696), .CLK(clk), .Q(ram[1259]) );
  DFFPOSX1 ram_reg_78__10_ ( .D(n5695), .CLK(clk), .Q(ram[1258]) );
  DFFPOSX1 ram_reg_78__9_ ( .D(n5694), .CLK(clk), .Q(ram[1257]) );
  DFFPOSX1 ram_reg_78__8_ ( .D(n5693), .CLK(clk), .Q(ram[1256]) );
  DFFPOSX1 ram_reg_78__7_ ( .D(n5692), .CLK(clk), .Q(ram[1255]) );
  DFFPOSX1 ram_reg_78__6_ ( .D(n5691), .CLK(clk), .Q(ram[1254]) );
  DFFPOSX1 ram_reg_78__5_ ( .D(n5690), .CLK(clk), .Q(ram[1253]) );
  DFFPOSX1 ram_reg_78__4_ ( .D(n5689), .CLK(clk), .Q(ram[1252]) );
  DFFPOSX1 ram_reg_78__3_ ( .D(n5688), .CLK(clk), .Q(ram[1251]) );
  DFFPOSX1 ram_reg_78__2_ ( .D(n5687), .CLK(clk), .Q(ram[1250]) );
  DFFPOSX1 ram_reg_78__1_ ( .D(n5686), .CLK(clk), .Q(ram[1249]) );
  DFFPOSX1 ram_reg_78__0_ ( .D(n5685), .CLK(clk), .Q(ram[1248]) );
  DFFPOSX1 ram_reg_77__15_ ( .D(n5684), .CLK(clk), .Q(ram[1247]) );
  DFFPOSX1 ram_reg_77__14_ ( .D(n5683), .CLK(clk), .Q(ram[1246]) );
  DFFPOSX1 ram_reg_77__13_ ( .D(n5682), .CLK(clk), .Q(ram[1245]) );
  DFFPOSX1 ram_reg_77__12_ ( .D(n5681), .CLK(clk), .Q(ram[1244]) );
  DFFPOSX1 ram_reg_77__11_ ( .D(n5680), .CLK(clk), .Q(ram[1243]) );
  DFFPOSX1 ram_reg_77__10_ ( .D(n5679), .CLK(clk), .Q(ram[1242]) );
  DFFPOSX1 ram_reg_77__9_ ( .D(n5678), .CLK(clk), .Q(ram[1241]) );
  DFFPOSX1 ram_reg_77__8_ ( .D(n5677), .CLK(clk), .Q(ram[1240]) );
  DFFPOSX1 ram_reg_77__7_ ( .D(n5676), .CLK(clk), .Q(ram[1239]) );
  DFFPOSX1 ram_reg_77__6_ ( .D(n5675), .CLK(clk), .Q(ram[1238]) );
  DFFPOSX1 ram_reg_77__5_ ( .D(n5674), .CLK(clk), .Q(ram[1237]) );
  DFFPOSX1 ram_reg_77__4_ ( .D(n5673), .CLK(clk), .Q(ram[1236]) );
  DFFPOSX1 ram_reg_77__3_ ( .D(n5672), .CLK(clk), .Q(ram[1235]) );
  DFFPOSX1 ram_reg_77__2_ ( .D(n5671), .CLK(clk), .Q(ram[1234]) );
  DFFPOSX1 ram_reg_77__1_ ( .D(n5670), .CLK(clk), .Q(ram[1233]) );
  DFFPOSX1 ram_reg_77__0_ ( .D(n5669), .CLK(clk), .Q(ram[1232]) );
  DFFPOSX1 ram_reg_76__15_ ( .D(n5668), .CLK(clk), .Q(ram[1231]) );
  DFFPOSX1 ram_reg_76__14_ ( .D(n5667), .CLK(clk), .Q(ram[1230]) );
  DFFPOSX1 ram_reg_76__13_ ( .D(n5666), .CLK(clk), .Q(ram[1229]) );
  DFFPOSX1 ram_reg_76__12_ ( .D(n5665), .CLK(clk), .Q(ram[1228]) );
  DFFPOSX1 ram_reg_76__11_ ( .D(n5664), .CLK(clk), .Q(ram[1227]) );
  DFFPOSX1 ram_reg_76__10_ ( .D(n5663), .CLK(clk), .Q(ram[1226]) );
  DFFPOSX1 ram_reg_76__9_ ( .D(n5662), .CLK(clk), .Q(ram[1225]) );
  DFFPOSX1 ram_reg_76__8_ ( .D(n5661), .CLK(clk), .Q(ram[1224]) );
  DFFPOSX1 ram_reg_76__7_ ( .D(n5660), .CLK(clk), .Q(ram[1223]) );
  DFFPOSX1 ram_reg_76__6_ ( .D(n5659), .CLK(clk), .Q(ram[1222]) );
  DFFPOSX1 ram_reg_76__5_ ( .D(n5658), .CLK(clk), .Q(ram[1221]) );
  DFFPOSX1 ram_reg_76__4_ ( .D(n5657), .CLK(clk), .Q(ram[1220]) );
  DFFPOSX1 ram_reg_76__3_ ( .D(n5656), .CLK(clk), .Q(ram[1219]) );
  DFFPOSX1 ram_reg_76__2_ ( .D(n5655), .CLK(clk), .Q(ram[1218]) );
  DFFPOSX1 ram_reg_76__1_ ( .D(n5654), .CLK(clk), .Q(ram[1217]) );
  DFFPOSX1 ram_reg_76__0_ ( .D(n5653), .CLK(clk), .Q(ram[1216]) );
  DFFPOSX1 ram_reg_75__15_ ( .D(n5652), .CLK(clk), .Q(ram[1215]) );
  DFFPOSX1 ram_reg_75__14_ ( .D(n5651), .CLK(clk), .Q(ram[1214]) );
  DFFPOSX1 ram_reg_75__13_ ( .D(n5650), .CLK(clk), .Q(ram[1213]) );
  DFFPOSX1 ram_reg_75__12_ ( .D(n5649), .CLK(clk), .Q(ram[1212]) );
  DFFPOSX1 ram_reg_75__11_ ( .D(n5648), .CLK(clk), .Q(ram[1211]) );
  DFFPOSX1 ram_reg_75__10_ ( .D(n5647), .CLK(clk), .Q(ram[1210]) );
  DFFPOSX1 ram_reg_75__9_ ( .D(n5646), .CLK(clk), .Q(ram[1209]) );
  DFFPOSX1 ram_reg_75__8_ ( .D(n5645), .CLK(clk), .Q(ram[1208]) );
  DFFPOSX1 ram_reg_75__7_ ( .D(n5644), .CLK(clk), .Q(ram[1207]) );
  DFFPOSX1 ram_reg_75__6_ ( .D(n5643), .CLK(clk), .Q(ram[1206]) );
  DFFPOSX1 ram_reg_75__5_ ( .D(n5642), .CLK(clk), .Q(ram[1205]) );
  DFFPOSX1 ram_reg_75__4_ ( .D(n5641), .CLK(clk), .Q(ram[1204]) );
  DFFPOSX1 ram_reg_75__3_ ( .D(n5640), .CLK(clk), .Q(ram[1203]) );
  DFFPOSX1 ram_reg_75__2_ ( .D(n5639), .CLK(clk), .Q(ram[1202]) );
  DFFPOSX1 ram_reg_75__1_ ( .D(n5638), .CLK(clk), .Q(ram[1201]) );
  DFFPOSX1 ram_reg_75__0_ ( .D(n5637), .CLK(clk), .Q(ram[1200]) );
  DFFPOSX1 ram_reg_74__15_ ( .D(n5636), .CLK(clk), .Q(ram[1199]) );
  DFFPOSX1 ram_reg_74__14_ ( .D(n5635), .CLK(clk), .Q(ram[1198]) );
  DFFPOSX1 ram_reg_74__13_ ( .D(n5634), .CLK(clk), .Q(ram[1197]) );
  DFFPOSX1 ram_reg_74__12_ ( .D(n5633), .CLK(clk), .Q(ram[1196]) );
  DFFPOSX1 ram_reg_74__11_ ( .D(n5632), .CLK(clk), .Q(ram[1195]) );
  DFFPOSX1 ram_reg_74__10_ ( .D(n5631), .CLK(clk), .Q(ram[1194]) );
  DFFPOSX1 ram_reg_74__9_ ( .D(n5630), .CLK(clk), .Q(ram[1193]) );
  DFFPOSX1 ram_reg_74__8_ ( .D(n5629), .CLK(clk), .Q(ram[1192]) );
  DFFPOSX1 ram_reg_74__7_ ( .D(n5628), .CLK(clk), .Q(ram[1191]) );
  DFFPOSX1 ram_reg_74__6_ ( .D(n5627), .CLK(clk), .Q(ram[1190]) );
  DFFPOSX1 ram_reg_74__5_ ( .D(n5626), .CLK(clk), .Q(ram[1189]) );
  DFFPOSX1 ram_reg_74__4_ ( .D(n5625), .CLK(clk), .Q(ram[1188]) );
  DFFPOSX1 ram_reg_74__3_ ( .D(n5624), .CLK(clk), .Q(ram[1187]) );
  DFFPOSX1 ram_reg_74__2_ ( .D(n5623), .CLK(clk), .Q(ram[1186]) );
  DFFPOSX1 ram_reg_74__1_ ( .D(n5622), .CLK(clk), .Q(ram[1185]) );
  DFFPOSX1 ram_reg_74__0_ ( .D(n5621), .CLK(clk), .Q(ram[1184]) );
  DFFPOSX1 ram_reg_73__15_ ( .D(n5620), .CLK(clk), .Q(ram[1183]) );
  DFFPOSX1 ram_reg_73__14_ ( .D(n5619), .CLK(clk), .Q(ram[1182]) );
  DFFPOSX1 ram_reg_73__13_ ( .D(n5618), .CLK(clk), .Q(ram[1181]) );
  DFFPOSX1 ram_reg_73__12_ ( .D(n5617), .CLK(clk), .Q(ram[1180]) );
  DFFPOSX1 ram_reg_73__11_ ( .D(n5616), .CLK(clk), .Q(ram[1179]) );
  DFFPOSX1 ram_reg_73__10_ ( .D(n5615), .CLK(clk), .Q(ram[1178]) );
  DFFPOSX1 ram_reg_73__9_ ( .D(n5614), .CLK(clk), .Q(ram[1177]) );
  DFFPOSX1 ram_reg_73__8_ ( .D(n5613), .CLK(clk), .Q(ram[1176]) );
  DFFPOSX1 ram_reg_73__7_ ( .D(n5612), .CLK(clk), .Q(ram[1175]) );
  DFFPOSX1 ram_reg_73__6_ ( .D(n5611), .CLK(clk), .Q(ram[1174]) );
  DFFPOSX1 ram_reg_73__5_ ( .D(n5610), .CLK(clk), .Q(ram[1173]) );
  DFFPOSX1 ram_reg_73__4_ ( .D(n5609), .CLK(clk), .Q(ram[1172]) );
  DFFPOSX1 ram_reg_73__3_ ( .D(n5608), .CLK(clk), .Q(ram[1171]) );
  DFFPOSX1 ram_reg_73__2_ ( .D(n5607), .CLK(clk), .Q(ram[1170]) );
  DFFPOSX1 ram_reg_73__1_ ( .D(n5606), .CLK(clk), .Q(ram[1169]) );
  DFFPOSX1 ram_reg_73__0_ ( .D(n5605), .CLK(clk), .Q(ram[1168]) );
  DFFPOSX1 ram_reg_72__15_ ( .D(n5604), .CLK(clk), .Q(ram[1167]) );
  DFFPOSX1 ram_reg_72__14_ ( .D(n5603), .CLK(clk), .Q(ram[1166]) );
  DFFPOSX1 ram_reg_72__13_ ( .D(n5602), .CLK(clk), .Q(ram[1165]) );
  DFFPOSX1 ram_reg_72__12_ ( .D(n5601), .CLK(clk), .Q(ram[1164]) );
  DFFPOSX1 ram_reg_72__11_ ( .D(n5600), .CLK(clk), .Q(ram[1163]) );
  DFFPOSX1 ram_reg_72__10_ ( .D(n5599), .CLK(clk), .Q(ram[1162]) );
  DFFPOSX1 ram_reg_72__9_ ( .D(n5598), .CLK(clk), .Q(ram[1161]) );
  DFFPOSX1 ram_reg_72__8_ ( .D(n5597), .CLK(clk), .Q(ram[1160]) );
  DFFPOSX1 ram_reg_72__7_ ( .D(n5596), .CLK(clk), .Q(ram[1159]) );
  DFFPOSX1 ram_reg_72__6_ ( .D(n5595), .CLK(clk), .Q(ram[1158]) );
  DFFPOSX1 ram_reg_72__5_ ( .D(n5594), .CLK(clk), .Q(ram[1157]) );
  DFFPOSX1 ram_reg_72__4_ ( .D(n5593), .CLK(clk), .Q(ram[1156]) );
  DFFPOSX1 ram_reg_72__3_ ( .D(n5592), .CLK(clk), .Q(ram[1155]) );
  DFFPOSX1 ram_reg_72__2_ ( .D(n5591), .CLK(clk), .Q(ram[1154]) );
  DFFPOSX1 ram_reg_72__1_ ( .D(n5590), .CLK(clk), .Q(ram[1153]) );
  DFFPOSX1 ram_reg_72__0_ ( .D(n5589), .CLK(clk), .Q(ram[1152]) );
  DFFPOSX1 ram_reg_71__15_ ( .D(n5588), .CLK(clk), .Q(ram[1151]) );
  DFFPOSX1 ram_reg_71__14_ ( .D(n5587), .CLK(clk), .Q(ram[1150]) );
  DFFPOSX1 ram_reg_71__13_ ( .D(n5586), .CLK(clk), .Q(ram[1149]) );
  DFFPOSX1 ram_reg_71__12_ ( .D(n5585), .CLK(clk), .Q(ram[1148]) );
  DFFPOSX1 ram_reg_71__11_ ( .D(n5584), .CLK(clk), .Q(ram[1147]) );
  DFFPOSX1 ram_reg_71__10_ ( .D(n5583), .CLK(clk), .Q(ram[1146]) );
  DFFPOSX1 ram_reg_71__9_ ( .D(n5582), .CLK(clk), .Q(ram[1145]) );
  DFFPOSX1 ram_reg_71__8_ ( .D(n5581), .CLK(clk), .Q(ram[1144]) );
  DFFPOSX1 ram_reg_71__7_ ( .D(n5580), .CLK(clk), .Q(ram[1143]) );
  DFFPOSX1 ram_reg_71__6_ ( .D(n5579), .CLK(clk), .Q(ram[1142]) );
  DFFPOSX1 ram_reg_71__5_ ( .D(n5578), .CLK(clk), .Q(ram[1141]) );
  DFFPOSX1 ram_reg_71__4_ ( .D(n5577), .CLK(clk), .Q(ram[1140]) );
  DFFPOSX1 ram_reg_71__3_ ( .D(n5576), .CLK(clk), .Q(ram[1139]) );
  DFFPOSX1 ram_reg_71__2_ ( .D(n5575), .CLK(clk), .Q(ram[1138]) );
  DFFPOSX1 ram_reg_71__1_ ( .D(n5574), .CLK(clk), .Q(ram[1137]) );
  DFFPOSX1 ram_reg_71__0_ ( .D(n5573), .CLK(clk), .Q(ram[1136]) );
  DFFPOSX1 ram_reg_70__15_ ( .D(n5572), .CLK(clk), .Q(ram[1135]) );
  DFFPOSX1 ram_reg_70__14_ ( .D(n5571), .CLK(clk), .Q(ram[1134]) );
  DFFPOSX1 ram_reg_70__13_ ( .D(n5570), .CLK(clk), .Q(ram[1133]) );
  DFFPOSX1 ram_reg_70__12_ ( .D(n5569), .CLK(clk), .Q(ram[1132]) );
  DFFPOSX1 ram_reg_70__11_ ( .D(n5568), .CLK(clk), .Q(ram[1131]) );
  DFFPOSX1 ram_reg_70__10_ ( .D(n5567), .CLK(clk), .Q(ram[1130]) );
  DFFPOSX1 ram_reg_70__9_ ( .D(n5566), .CLK(clk), .Q(ram[1129]) );
  DFFPOSX1 ram_reg_70__8_ ( .D(n5565), .CLK(clk), .Q(ram[1128]) );
  DFFPOSX1 ram_reg_70__7_ ( .D(n5564), .CLK(clk), .Q(ram[1127]) );
  DFFPOSX1 ram_reg_70__6_ ( .D(n5563), .CLK(clk), .Q(ram[1126]) );
  DFFPOSX1 ram_reg_70__5_ ( .D(n5562), .CLK(clk), .Q(ram[1125]) );
  DFFPOSX1 ram_reg_70__4_ ( .D(n5561), .CLK(clk), .Q(ram[1124]) );
  DFFPOSX1 ram_reg_70__3_ ( .D(n5560), .CLK(clk), .Q(ram[1123]) );
  DFFPOSX1 ram_reg_70__2_ ( .D(n5559), .CLK(clk), .Q(ram[1122]) );
  DFFPOSX1 ram_reg_70__1_ ( .D(n5558), .CLK(clk), .Q(ram[1121]) );
  DFFPOSX1 ram_reg_70__0_ ( .D(n5557), .CLK(clk), .Q(ram[1120]) );
  DFFPOSX1 ram_reg_69__15_ ( .D(n5556), .CLK(clk), .Q(ram[1119]) );
  DFFPOSX1 ram_reg_69__14_ ( .D(n5555), .CLK(clk), .Q(ram[1118]) );
  DFFPOSX1 ram_reg_69__13_ ( .D(n5554), .CLK(clk), .Q(ram[1117]) );
  DFFPOSX1 ram_reg_69__12_ ( .D(n5553), .CLK(clk), .Q(ram[1116]) );
  DFFPOSX1 ram_reg_69__11_ ( .D(n5552), .CLK(clk), .Q(ram[1115]) );
  DFFPOSX1 ram_reg_69__10_ ( .D(n5551), .CLK(clk), .Q(ram[1114]) );
  DFFPOSX1 ram_reg_69__9_ ( .D(n5550), .CLK(clk), .Q(ram[1113]) );
  DFFPOSX1 ram_reg_69__8_ ( .D(n5549), .CLK(clk), .Q(ram[1112]) );
  DFFPOSX1 ram_reg_69__7_ ( .D(n5548), .CLK(clk), .Q(ram[1111]) );
  DFFPOSX1 ram_reg_69__6_ ( .D(n5547), .CLK(clk), .Q(ram[1110]) );
  DFFPOSX1 ram_reg_69__5_ ( .D(n5546), .CLK(clk), .Q(ram[1109]) );
  DFFPOSX1 ram_reg_69__4_ ( .D(n5545), .CLK(clk), .Q(ram[1108]) );
  DFFPOSX1 ram_reg_69__3_ ( .D(n5544), .CLK(clk), .Q(ram[1107]) );
  DFFPOSX1 ram_reg_69__2_ ( .D(n5543), .CLK(clk), .Q(ram[1106]) );
  DFFPOSX1 ram_reg_69__1_ ( .D(n5542), .CLK(clk), .Q(ram[1105]) );
  DFFPOSX1 ram_reg_69__0_ ( .D(n5541), .CLK(clk), .Q(ram[1104]) );
  DFFPOSX1 ram_reg_68__15_ ( .D(n5540), .CLK(clk), .Q(ram[1103]) );
  DFFPOSX1 ram_reg_68__14_ ( .D(n5539), .CLK(clk), .Q(ram[1102]) );
  DFFPOSX1 ram_reg_68__13_ ( .D(n5538), .CLK(clk), .Q(ram[1101]) );
  DFFPOSX1 ram_reg_68__12_ ( .D(n5537), .CLK(clk), .Q(ram[1100]) );
  DFFPOSX1 ram_reg_68__11_ ( .D(n5536), .CLK(clk), .Q(ram[1099]) );
  DFFPOSX1 ram_reg_68__10_ ( .D(n5535), .CLK(clk), .Q(ram[1098]) );
  DFFPOSX1 ram_reg_68__9_ ( .D(n5534), .CLK(clk), .Q(ram[1097]) );
  DFFPOSX1 ram_reg_68__8_ ( .D(n5533), .CLK(clk), .Q(ram[1096]) );
  DFFPOSX1 ram_reg_68__7_ ( .D(n5532), .CLK(clk), .Q(ram[1095]) );
  DFFPOSX1 ram_reg_68__6_ ( .D(n5531), .CLK(clk), .Q(ram[1094]) );
  DFFPOSX1 ram_reg_68__5_ ( .D(n5530), .CLK(clk), .Q(ram[1093]) );
  DFFPOSX1 ram_reg_68__4_ ( .D(n5529), .CLK(clk), .Q(ram[1092]) );
  DFFPOSX1 ram_reg_68__3_ ( .D(n5528), .CLK(clk), .Q(ram[1091]) );
  DFFPOSX1 ram_reg_68__2_ ( .D(n5527), .CLK(clk), .Q(ram[1090]) );
  DFFPOSX1 ram_reg_68__1_ ( .D(n5526), .CLK(clk), .Q(ram[1089]) );
  DFFPOSX1 ram_reg_68__0_ ( .D(n5525), .CLK(clk), .Q(ram[1088]) );
  DFFPOSX1 ram_reg_67__15_ ( .D(n5524), .CLK(clk), .Q(ram[1087]) );
  DFFPOSX1 ram_reg_67__14_ ( .D(n5523), .CLK(clk), .Q(ram[1086]) );
  DFFPOSX1 ram_reg_67__13_ ( .D(n5522), .CLK(clk), .Q(ram[1085]) );
  DFFPOSX1 ram_reg_67__12_ ( .D(n5521), .CLK(clk), .Q(ram[1084]) );
  DFFPOSX1 ram_reg_67__11_ ( .D(n5520), .CLK(clk), .Q(ram[1083]) );
  DFFPOSX1 ram_reg_67__10_ ( .D(n5519), .CLK(clk), .Q(ram[1082]) );
  DFFPOSX1 ram_reg_67__9_ ( .D(n5518), .CLK(clk), .Q(ram[1081]) );
  DFFPOSX1 ram_reg_67__8_ ( .D(n5517), .CLK(clk), .Q(ram[1080]) );
  DFFPOSX1 ram_reg_67__7_ ( .D(n5516), .CLK(clk), .Q(ram[1079]) );
  DFFPOSX1 ram_reg_67__6_ ( .D(n5515), .CLK(clk), .Q(ram[1078]) );
  DFFPOSX1 ram_reg_67__5_ ( .D(n5514), .CLK(clk), .Q(ram[1077]) );
  DFFPOSX1 ram_reg_67__4_ ( .D(n5513), .CLK(clk), .Q(ram[1076]) );
  DFFPOSX1 ram_reg_67__3_ ( .D(n5512), .CLK(clk), .Q(ram[1075]) );
  DFFPOSX1 ram_reg_67__2_ ( .D(n5511), .CLK(clk), .Q(ram[1074]) );
  DFFPOSX1 ram_reg_67__1_ ( .D(n5510), .CLK(clk), .Q(ram[1073]) );
  DFFPOSX1 ram_reg_67__0_ ( .D(n5509), .CLK(clk), .Q(ram[1072]) );
  DFFPOSX1 ram_reg_66__15_ ( .D(n5508), .CLK(clk), .Q(ram[1071]) );
  DFFPOSX1 ram_reg_66__14_ ( .D(n5507), .CLK(clk), .Q(ram[1070]) );
  DFFPOSX1 ram_reg_66__13_ ( .D(n5506), .CLK(clk), .Q(ram[1069]) );
  DFFPOSX1 ram_reg_66__12_ ( .D(n5505), .CLK(clk), .Q(ram[1068]) );
  DFFPOSX1 ram_reg_66__11_ ( .D(n5504), .CLK(clk), .Q(ram[1067]) );
  DFFPOSX1 ram_reg_66__10_ ( .D(n5503), .CLK(clk), .Q(ram[1066]) );
  DFFPOSX1 ram_reg_66__9_ ( .D(n5502), .CLK(clk), .Q(ram[1065]) );
  DFFPOSX1 ram_reg_66__8_ ( .D(n5501), .CLK(clk), .Q(ram[1064]) );
  DFFPOSX1 ram_reg_66__7_ ( .D(n5500), .CLK(clk), .Q(ram[1063]) );
  DFFPOSX1 ram_reg_66__6_ ( .D(n5499), .CLK(clk), .Q(ram[1062]) );
  DFFPOSX1 ram_reg_66__5_ ( .D(n5498), .CLK(clk), .Q(ram[1061]) );
  DFFPOSX1 ram_reg_66__4_ ( .D(n5497), .CLK(clk), .Q(ram[1060]) );
  DFFPOSX1 ram_reg_66__3_ ( .D(n5496), .CLK(clk), .Q(ram[1059]) );
  DFFPOSX1 ram_reg_66__2_ ( .D(n5495), .CLK(clk), .Q(ram[1058]) );
  DFFPOSX1 ram_reg_66__1_ ( .D(n5494), .CLK(clk), .Q(ram[1057]) );
  DFFPOSX1 ram_reg_66__0_ ( .D(n5493), .CLK(clk), .Q(ram[1056]) );
  DFFPOSX1 ram_reg_65__15_ ( .D(n5492), .CLK(clk), .Q(ram[1055]) );
  DFFPOSX1 ram_reg_65__14_ ( .D(n5491), .CLK(clk), .Q(ram[1054]) );
  DFFPOSX1 ram_reg_65__13_ ( .D(n5490), .CLK(clk), .Q(ram[1053]) );
  DFFPOSX1 ram_reg_65__12_ ( .D(n5489), .CLK(clk), .Q(ram[1052]) );
  DFFPOSX1 ram_reg_65__11_ ( .D(n5488), .CLK(clk), .Q(ram[1051]) );
  DFFPOSX1 ram_reg_65__10_ ( .D(n5487), .CLK(clk), .Q(ram[1050]) );
  DFFPOSX1 ram_reg_65__9_ ( .D(n5486), .CLK(clk), .Q(ram[1049]) );
  DFFPOSX1 ram_reg_65__8_ ( .D(n5485), .CLK(clk), .Q(ram[1048]) );
  DFFPOSX1 ram_reg_65__7_ ( .D(n5484), .CLK(clk), .Q(ram[1047]) );
  DFFPOSX1 ram_reg_65__6_ ( .D(n5483), .CLK(clk), .Q(ram[1046]) );
  DFFPOSX1 ram_reg_65__5_ ( .D(n5482), .CLK(clk), .Q(ram[1045]) );
  DFFPOSX1 ram_reg_65__4_ ( .D(n5481), .CLK(clk), .Q(ram[1044]) );
  DFFPOSX1 ram_reg_65__3_ ( .D(n5480), .CLK(clk), .Q(ram[1043]) );
  DFFPOSX1 ram_reg_65__2_ ( .D(n5479), .CLK(clk), .Q(ram[1042]) );
  DFFPOSX1 ram_reg_65__1_ ( .D(n5478), .CLK(clk), .Q(ram[1041]) );
  DFFPOSX1 ram_reg_65__0_ ( .D(n5477), .CLK(clk), .Q(ram[1040]) );
  DFFPOSX1 ram_reg_64__15_ ( .D(n5476), .CLK(clk), .Q(ram[1039]) );
  DFFPOSX1 ram_reg_64__14_ ( .D(n5475), .CLK(clk), .Q(ram[1038]) );
  DFFPOSX1 ram_reg_64__13_ ( .D(n5474), .CLK(clk), .Q(ram[1037]) );
  DFFPOSX1 ram_reg_64__12_ ( .D(n5473), .CLK(clk), .Q(ram[1036]) );
  DFFPOSX1 ram_reg_64__11_ ( .D(n5472), .CLK(clk), .Q(ram[1035]) );
  DFFPOSX1 ram_reg_64__10_ ( .D(n5471), .CLK(clk), .Q(ram[1034]) );
  DFFPOSX1 ram_reg_64__9_ ( .D(n5470), .CLK(clk), .Q(ram[1033]) );
  DFFPOSX1 ram_reg_64__8_ ( .D(n5469), .CLK(clk), .Q(ram[1032]) );
  DFFPOSX1 ram_reg_64__7_ ( .D(n5468), .CLK(clk), .Q(ram[1031]) );
  DFFPOSX1 ram_reg_64__6_ ( .D(n5467), .CLK(clk), .Q(ram[1030]) );
  DFFPOSX1 ram_reg_64__5_ ( .D(n5466), .CLK(clk), .Q(ram[1029]) );
  DFFPOSX1 ram_reg_64__4_ ( .D(n5465), .CLK(clk), .Q(ram[1028]) );
  DFFPOSX1 ram_reg_64__3_ ( .D(n5464), .CLK(clk), .Q(ram[1027]) );
  DFFPOSX1 ram_reg_64__2_ ( .D(n5463), .CLK(clk), .Q(ram[1026]) );
  DFFPOSX1 ram_reg_64__1_ ( .D(n5462), .CLK(clk), .Q(ram[1025]) );
  DFFPOSX1 ram_reg_64__0_ ( .D(n5461), .CLK(clk), .Q(ram[1024]) );
  DFFPOSX1 ram_reg_63__15_ ( .D(n5460), .CLK(clk), .Q(ram[1023]) );
  DFFPOSX1 ram_reg_63__14_ ( .D(n5459), .CLK(clk), .Q(ram[1022]) );
  DFFPOSX1 ram_reg_63__13_ ( .D(n5458), .CLK(clk), .Q(ram[1021]) );
  DFFPOSX1 ram_reg_63__12_ ( .D(n5457), .CLK(clk), .Q(ram[1020]) );
  DFFPOSX1 ram_reg_63__11_ ( .D(n5456), .CLK(clk), .Q(ram[1019]) );
  DFFPOSX1 ram_reg_63__10_ ( .D(n5455), .CLK(clk), .Q(ram[1018]) );
  DFFPOSX1 ram_reg_63__9_ ( .D(n5454), .CLK(clk), .Q(ram[1017]) );
  DFFPOSX1 ram_reg_63__8_ ( .D(n5453), .CLK(clk), .Q(ram[1016]) );
  DFFPOSX1 ram_reg_63__7_ ( .D(n5452), .CLK(clk), .Q(ram[1015]) );
  DFFPOSX1 ram_reg_63__6_ ( .D(n5451), .CLK(clk), .Q(ram[1014]) );
  DFFPOSX1 ram_reg_63__5_ ( .D(n5450), .CLK(clk), .Q(ram[1013]) );
  DFFPOSX1 ram_reg_63__4_ ( .D(n5449), .CLK(clk), .Q(ram[1012]) );
  DFFPOSX1 ram_reg_63__3_ ( .D(n5448), .CLK(clk), .Q(ram[1011]) );
  DFFPOSX1 ram_reg_63__2_ ( .D(n5447), .CLK(clk), .Q(ram[1010]) );
  DFFPOSX1 ram_reg_63__1_ ( .D(n5446), .CLK(clk), .Q(ram[1009]) );
  DFFPOSX1 ram_reg_63__0_ ( .D(n5445), .CLK(clk), .Q(ram[1008]) );
  DFFPOSX1 ram_reg_62__15_ ( .D(n5444), .CLK(clk), .Q(ram[1007]) );
  DFFPOSX1 ram_reg_62__14_ ( .D(n5443), .CLK(clk), .Q(ram[1006]) );
  DFFPOSX1 ram_reg_62__13_ ( .D(n5442), .CLK(clk), .Q(ram[1005]) );
  DFFPOSX1 ram_reg_62__12_ ( .D(n5441), .CLK(clk), .Q(ram[1004]) );
  DFFPOSX1 ram_reg_62__11_ ( .D(n5440), .CLK(clk), .Q(ram[1003]) );
  DFFPOSX1 ram_reg_62__10_ ( .D(n5439), .CLK(clk), .Q(ram[1002]) );
  DFFPOSX1 ram_reg_62__9_ ( .D(n5438), .CLK(clk), .Q(ram[1001]) );
  DFFPOSX1 ram_reg_62__8_ ( .D(n5437), .CLK(clk), .Q(ram[1000]) );
  DFFPOSX1 ram_reg_62__7_ ( .D(n5436), .CLK(clk), .Q(ram[999]) );
  DFFPOSX1 ram_reg_62__6_ ( .D(n5435), .CLK(clk), .Q(ram[998]) );
  DFFPOSX1 ram_reg_62__5_ ( .D(n5434), .CLK(clk), .Q(ram[997]) );
  DFFPOSX1 ram_reg_62__4_ ( .D(n5433), .CLK(clk), .Q(ram[996]) );
  DFFPOSX1 ram_reg_62__3_ ( .D(n5432), .CLK(clk), .Q(ram[995]) );
  DFFPOSX1 ram_reg_62__2_ ( .D(n5431), .CLK(clk), .Q(ram[994]) );
  DFFPOSX1 ram_reg_62__1_ ( .D(n5430), .CLK(clk), .Q(ram[993]) );
  DFFPOSX1 ram_reg_62__0_ ( .D(n5429), .CLK(clk), .Q(ram[992]) );
  DFFPOSX1 ram_reg_61__15_ ( .D(n5428), .CLK(clk), .Q(ram[991]) );
  DFFPOSX1 ram_reg_61__14_ ( .D(n5427), .CLK(clk), .Q(ram[990]) );
  DFFPOSX1 ram_reg_61__13_ ( .D(n5426), .CLK(clk), .Q(ram[989]) );
  DFFPOSX1 ram_reg_61__12_ ( .D(n5425), .CLK(clk), .Q(ram[988]) );
  DFFPOSX1 ram_reg_61__11_ ( .D(n5424), .CLK(clk), .Q(ram[987]) );
  DFFPOSX1 ram_reg_61__10_ ( .D(n5423), .CLK(clk), .Q(ram[986]) );
  DFFPOSX1 ram_reg_61__9_ ( .D(n5422), .CLK(clk), .Q(ram[985]) );
  DFFPOSX1 ram_reg_61__8_ ( .D(n5421), .CLK(clk), .Q(ram[984]) );
  DFFPOSX1 ram_reg_61__7_ ( .D(n5420), .CLK(clk), .Q(ram[983]) );
  DFFPOSX1 ram_reg_61__6_ ( .D(n5419), .CLK(clk), .Q(ram[982]) );
  DFFPOSX1 ram_reg_61__5_ ( .D(n5418), .CLK(clk), .Q(ram[981]) );
  DFFPOSX1 ram_reg_61__4_ ( .D(n5417), .CLK(clk), .Q(ram[980]) );
  DFFPOSX1 ram_reg_61__3_ ( .D(n5416), .CLK(clk), .Q(ram[979]) );
  DFFPOSX1 ram_reg_61__2_ ( .D(n5415), .CLK(clk), .Q(ram[978]) );
  DFFPOSX1 ram_reg_61__1_ ( .D(n5414), .CLK(clk), .Q(ram[977]) );
  DFFPOSX1 ram_reg_61__0_ ( .D(n5413), .CLK(clk), .Q(ram[976]) );
  DFFPOSX1 ram_reg_60__15_ ( .D(n5412), .CLK(clk), .Q(ram[975]) );
  DFFPOSX1 ram_reg_60__14_ ( .D(n5411), .CLK(clk), .Q(ram[974]) );
  DFFPOSX1 ram_reg_60__13_ ( .D(n5410), .CLK(clk), .Q(ram[973]) );
  DFFPOSX1 ram_reg_60__12_ ( .D(n5409), .CLK(clk), .Q(ram[972]) );
  DFFPOSX1 ram_reg_60__11_ ( .D(n5408), .CLK(clk), .Q(ram[971]) );
  DFFPOSX1 ram_reg_60__10_ ( .D(n5407), .CLK(clk), .Q(ram[970]) );
  DFFPOSX1 ram_reg_60__9_ ( .D(n5406), .CLK(clk), .Q(ram[969]) );
  DFFPOSX1 ram_reg_60__8_ ( .D(n5405), .CLK(clk), .Q(ram[968]) );
  DFFPOSX1 ram_reg_60__7_ ( .D(n5404), .CLK(clk), .Q(ram[967]) );
  DFFPOSX1 ram_reg_60__6_ ( .D(n5403), .CLK(clk), .Q(ram[966]) );
  DFFPOSX1 ram_reg_60__5_ ( .D(n5402), .CLK(clk), .Q(ram[965]) );
  DFFPOSX1 ram_reg_60__4_ ( .D(n5401), .CLK(clk), .Q(ram[964]) );
  DFFPOSX1 ram_reg_60__3_ ( .D(n5400), .CLK(clk), .Q(ram[963]) );
  DFFPOSX1 ram_reg_60__2_ ( .D(n5399), .CLK(clk), .Q(ram[962]) );
  DFFPOSX1 ram_reg_60__1_ ( .D(n5398), .CLK(clk), .Q(ram[961]) );
  DFFPOSX1 ram_reg_60__0_ ( .D(n5397), .CLK(clk), .Q(ram[960]) );
  DFFPOSX1 ram_reg_59__15_ ( .D(n5396), .CLK(clk), .Q(ram[959]) );
  DFFPOSX1 ram_reg_59__14_ ( .D(n5395), .CLK(clk), .Q(ram[958]) );
  DFFPOSX1 ram_reg_59__13_ ( .D(n5394), .CLK(clk), .Q(ram[957]) );
  DFFPOSX1 ram_reg_59__12_ ( .D(n5393), .CLK(clk), .Q(ram[956]) );
  DFFPOSX1 ram_reg_59__11_ ( .D(n5392), .CLK(clk), .Q(ram[955]) );
  DFFPOSX1 ram_reg_59__10_ ( .D(n5391), .CLK(clk), .Q(ram[954]) );
  DFFPOSX1 ram_reg_59__9_ ( .D(n5390), .CLK(clk), .Q(ram[953]) );
  DFFPOSX1 ram_reg_59__8_ ( .D(n5389), .CLK(clk), .Q(ram[952]) );
  DFFPOSX1 ram_reg_59__7_ ( .D(n5388), .CLK(clk), .Q(ram[951]) );
  DFFPOSX1 ram_reg_59__6_ ( .D(n5387), .CLK(clk), .Q(ram[950]) );
  DFFPOSX1 ram_reg_59__5_ ( .D(n5386), .CLK(clk), .Q(ram[949]) );
  DFFPOSX1 ram_reg_59__4_ ( .D(n5385), .CLK(clk), .Q(ram[948]) );
  DFFPOSX1 ram_reg_59__3_ ( .D(n5384), .CLK(clk), .Q(ram[947]) );
  DFFPOSX1 ram_reg_59__2_ ( .D(n5383), .CLK(clk), .Q(ram[946]) );
  DFFPOSX1 ram_reg_59__1_ ( .D(n5382), .CLK(clk), .Q(ram[945]) );
  DFFPOSX1 ram_reg_59__0_ ( .D(n5381), .CLK(clk), .Q(ram[944]) );
  DFFPOSX1 ram_reg_58__15_ ( .D(n5380), .CLK(clk), .Q(ram[943]) );
  DFFPOSX1 ram_reg_58__14_ ( .D(n5379), .CLK(clk), .Q(ram[942]) );
  DFFPOSX1 ram_reg_58__13_ ( .D(n5378), .CLK(clk), .Q(ram[941]) );
  DFFPOSX1 ram_reg_58__12_ ( .D(n5377), .CLK(clk), .Q(ram[940]) );
  DFFPOSX1 ram_reg_58__11_ ( .D(n5376), .CLK(clk), .Q(ram[939]) );
  DFFPOSX1 ram_reg_58__10_ ( .D(n5375), .CLK(clk), .Q(ram[938]) );
  DFFPOSX1 ram_reg_58__9_ ( .D(n5374), .CLK(clk), .Q(ram[937]) );
  DFFPOSX1 ram_reg_58__8_ ( .D(n5373), .CLK(clk), .Q(ram[936]) );
  DFFPOSX1 ram_reg_58__7_ ( .D(n5372), .CLK(clk), .Q(ram[935]) );
  DFFPOSX1 ram_reg_58__6_ ( .D(n5371), .CLK(clk), .Q(ram[934]) );
  DFFPOSX1 ram_reg_58__5_ ( .D(n5370), .CLK(clk), .Q(ram[933]) );
  DFFPOSX1 ram_reg_58__4_ ( .D(n5369), .CLK(clk), .Q(ram[932]) );
  DFFPOSX1 ram_reg_58__3_ ( .D(n5368), .CLK(clk), .Q(ram[931]) );
  DFFPOSX1 ram_reg_58__2_ ( .D(n5367), .CLK(clk), .Q(ram[930]) );
  DFFPOSX1 ram_reg_58__1_ ( .D(n5366), .CLK(clk), .Q(ram[929]) );
  DFFPOSX1 ram_reg_58__0_ ( .D(n5365), .CLK(clk), .Q(ram[928]) );
  DFFPOSX1 ram_reg_57__15_ ( .D(n5364), .CLK(clk), .Q(ram[927]) );
  DFFPOSX1 ram_reg_57__14_ ( .D(n5363), .CLK(clk), .Q(ram[926]) );
  DFFPOSX1 ram_reg_57__13_ ( .D(n5362), .CLK(clk), .Q(ram[925]) );
  DFFPOSX1 ram_reg_57__12_ ( .D(n5361), .CLK(clk), .Q(ram[924]) );
  DFFPOSX1 ram_reg_57__11_ ( .D(n5360), .CLK(clk), .Q(ram[923]) );
  DFFPOSX1 ram_reg_57__10_ ( .D(n5359), .CLK(clk), .Q(ram[922]) );
  DFFPOSX1 ram_reg_57__9_ ( .D(n5358), .CLK(clk), .Q(ram[921]) );
  DFFPOSX1 ram_reg_57__8_ ( .D(n5357), .CLK(clk), .Q(ram[920]) );
  DFFPOSX1 ram_reg_57__7_ ( .D(n5356), .CLK(clk), .Q(ram[919]) );
  DFFPOSX1 ram_reg_57__6_ ( .D(n5355), .CLK(clk), .Q(ram[918]) );
  DFFPOSX1 ram_reg_57__5_ ( .D(n5354), .CLK(clk), .Q(ram[917]) );
  DFFPOSX1 ram_reg_57__4_ ( .D(n5353), .CLK(clk), .Q(ram[916]) );
  DFFPOSX1 ram_reg_57__3_ ( .D(n5352), .CLK(clk), .Q(ram[915]) );
  DFFPOSX1 ram_reg_57__2_ ( .D(n5351), .CLK(clk), .Q(ram[914]) );
  DFFPOSX1 ram_reg_57__1_ ( .D(n5350), .CLK(clk), .Q(ram[913]) );
  DFFPOSX1 ram_reg_57__0_ ( .D(n5349), .CLK(clk), .Q(ram[912]) );
  DFFPOSX1 ram_reg_56__15_ ( .D(n5348), .CLK(clk), .Q(ram[911]) );
  DFFPOSX1 ram_reg_56__14_ ( .D(n5347), .CLK(clk), .Q(ram[910]) );
  DFFPOSX1 ram_reg_56__13_ ( .D(n5346), .CLK(clk), .Q(ram[909]) );
  DFFPOSX1 ram_reg_56__12_ ( .D(n5345), .CLK(clk), .Q(ram[908]) );
  DFFPOSX1 ram_reg_56__11_ ( .D(n5344), .CLK(clk), .Q(ram[907]) );
  DFFPOSX1 ram_reg_56__10_ ( .D(n5343), .CLK(clk), .Q(ram[906]) );
  DFFPOSX1 ram_reg_56__9_ ( .D(n5342), .CLK(clk), .Q(ram[905]) );
  DFFPOSX1 ram_reg_56__8_ ( .D(n5341), .CLK(clk), .Q(ram[904]) );
  DFFPOSX1 ram_reg_56__7_ ( .D(n5340), .CLK(clk), .Q(ram[903]) );
  DFFPOSX1 ram_reg_56__6_ ( .D(n5339), .CLK(clk), .Q(ram[902]) );
  DFFPOSX1 ram_reg_56__5_ ( .D(n5338), .CLK(clk), .Q(ram[901]) );
  DFFPOSX1 ram_reg_56__4_ ( .D(n5337), .CLK(clk), .Q(ram[900]) );
  DFFPOSX1 ram_reg_56__3_ ( .D(n5336), .CLK(clk), .Q(ram[899]) );
  DFFPOSX1 ram_reg_56__2_ ( .D(n5335), .CLK(clk), .Q(ram[898]) );
  DFFPOSX1 ram_reg_56__1_ ( .D(n5334), .CLK(clk), .Q(ram[897]) );
  DFFPOSX1 ram_reg_56__0_ ( .D(n5333), .CLK(clk), .Q(ram[896]) );
  DFFPOSX1 ram_reg_55__15_ ( .D(n5332), .CLK(clk), .Q(ram[895]) );
  DFFPOSX1 ram_reg_55__14_ ( .D(n5331), .CLK(clk), .Q(ram[894]) );
  DFFPOSX1 ram_reg_55__13_ ( .D(n5330), .CLK(clk), .Q(ram[893]) );
  DFFPOSX1 ram_reg_55__12_ ( .D(n5329), .CLK(clk), .Q(ram[892]) );
  DFFPOSX1 ram_reg_55__11_ ( .D(n5328), .CLK(clk), .Q(ram[891]) );
  DFFPOSX1 ram_reg_55__10_ ( .D(n5327), .CLK(clk), .Q(ram[890]) );
  DFFPOSX1 ram_reg_55__9_ ( .D(n5326), .CLK(clk), .Q(ram[889]) );
  DFFPOSX1 ram_reg_55__8_ ( .D(n5325), .CLK(clk), .Q(ram[888]) );
  DFFPOSX1 ram_reg_55__7_ ( .D(n5324), .CLK(clk), .Q(ram[887]) );
  DFFPOSX1 ram_reg_55__6_ ( .D(n5323), .CLK(clk), .Q(ram[886]) );
  DFFPOSX1 ram_reg_55__5_ ( .D(n5322), .CLK(clk), .Q(ram[885]) );
  DFFPOSX1 ram_reg_55__4_ ( .D(n5321), .CLK(clk), .Q(ram[884]) );
  DFFPOSX1 ram_reg_55__3_ ( .D(n5320), .CLK(clk), .Q(ram[883]) );
  DFFPOSX1 ram_reg_55__2_ ( .D(n5319), .CLK(clk), .Q(ram[882]) );
  DFFPOSX1 ram_reg_55__1_ ( .D(n5318), .CLK(clk), .Q(ram[881]) );
  DFFPOSX1 ram_reg_55__0_ ( .D(n5317), .CLK(clk), .Q(ram[880]) );
  DFFPOSX1 ram_reg_54__15_ ( .D(n5316), .CLK(clk), .Q(ram[879]) );
  DFFPOSX1 ram_reg_54__14_ ( .D(n5315), .CLK(clk), .Q(ram[878]) );
  DFFPOSX1 ram_reg_54__13_ ( .D(n5314), .CLK(clk), .Q(ram[877]) );
  DFFPOSX1 ram_reg_54__12_ ( .D(n5313), .CLK(clk), .Q(ram[876]) );
  DFFPOSX1 ram_reg_54__11_ ( .D(n5312), .CLK(clk), .Q(ram[875]) );
  DFFPOSX1 ram_reg_54__10_ ( .D(n5311), .CLK(clk), .Q(ram[874]) );
  DFFPOSX1 ram_reg_54__9_ ( .D(n5310), .CLK(clk), .Q(ram[873]) );
  DFFPOSX1 ram_reg_54__8_ ( .D(n5309), .CLK(clk), .Q(ram[872]) );
  DFFPOSX1 ram_reg_54__7_ ( .D(n5308), .CLK(clk), .Q(ram[871]) );
  DFFPOSX1 ram_reg_54__6_ ( .D(n5307), .CLK(clk), .Q(ram[870]) );
  DFFPOSX1 ram_reg_54__5_ ( .D(n5306), .CLK(clk), .Q(ram[869]) );
  DFFPOSX1 ram_reg_54__4_ ( .D(n5305), .CLK(clk), .Q(ram[868]) );
  DFFPOSX1 ram_reg_54__3_ ( .D(n5304), .CLK(clk), .Q(ram[867]) );
  DFFPOSX1 ram_reg_54__2_ ( .D(n5303), .CLK(clk), .Q(ram[866]) );
  DFFPOSX1 ram_reg_54__1_ ( .D(n5302), .CLK(clk), .Q(ram[865]) );
  DFFPOSX1 ram_reg_54__0_ ( .D(n5301), .CLK(clk), .Q(ram[864]) );
  DFFPOSX1 ram_reg_53__15_ ( .D(n5300), .CLK(clk), .Q(ram[863]) );
  DFFPOSX1 ram_reg_53__14_ ( .D(n5299), .CLK(clk), .Q(ram[862]) );
  DFFPOSX1 ram_reg_53__13_ ( .D(n5298), .CLK(clk), .Q(ram[861]) );
  DFFPOSX1 ram_reg_53__12_ ( .D(n5297), .CLK(clk), .Q(ram[860]) );
  DFFPOSX1 ram_reg_53__11_ ( .D(n5296), .CLK(clk), .Q(ram[859]) );
  DFFPOSX1 ram_reg_53__10_ ( .D(n5295), .CLK(clk), .Q(ram[858]) );
  DFFPOSX1 ram_reg_53__9_ ( .D(n5294), .CLK(clk), .Q(ram[857]) );
  DFFPOSX1 ram_reg_53__8_ ( .D(n5293), .CLK(clk), .Q(ram[856]) );
  DFFPOSX1 ram_reg_53__7_ ( .D(n5292), .CLK(clk), .Q(ram[855]) );
  DFFPOSX1 ram_reg_53__6_ ( .D(n5291), .CLK(clk), .Q(ram[854]) );
  DFFPOSX1 ram_reg_53__5_ ( .D(n5290), .CLK(clk), .Q(ram[853]) );
  DFFPOSX1 ram_reg_53__4_ ( .D(n5289), .CLK(clk), .Q(ram[852]) );
  DFFPOSX1 ram_reg_53__3_ ( .D(n5288), .CLK(clk), .Q(ram[851]) );
  DFFPOSX1 ram_reg_53__2_ ( .D(n5287), .CLK(clk), .Q(ram[850]) );
  DFFPOSX1 ram_reg_53__1_ ( .D(n5286), .CLK(clk), .Q(ram[849]) );
  DFFPOSX1 ram_reg_53__0_ ( .D(n5285), .CLK(clk), .Q(ram[848]) );
  DFFPOSX1 ram_reg_52__15_ ( .D(n5284), .CLK(clk), .Q(ram[847]) );
  DFFPOSX1 ram_reg_52__14_ ( .D(n5283), .CLK(clk), .Q(ram[846]) );
  DFFPOSX1 ram_reg_52__13_ ( .D(n5282), .CLK(clk), .Q(ram[845]) );
  DFFPOSX1 ram_reg_52__12_ ( .D(n5281), .CLK(clk), .Q(ram[844]) );
  DFFPOSX1 ram_reg_52__11_ ( .D(n5280), .CLK(clk), .Q(ram[843]) );
  DFFPOSX1 ram_reg_52__10_ ( .D(n5279), .CLK(clk), .Q(ram[842]) );
  DFFPOSX1 ram_reg_52__9_ ( .D(n5278), .CLK(clk), .Q(ram[841]) );
  DFFPOSX1 ram_reg_52__8_ ( .D(n5277), .CLK(clk), .Q(ram[840]) );
  DFFPOSX1 ram_reg_52__7_ ( .D(n5276), .CLK(clk), .Q(ram[839]) );
  DFFPOSX1 ram_reg_52__6_ ( .D(n5275), .CLK(clk), .Q(ram[838]) );
  DFFPOSX1 ram_reg_52__5_ ( .D(n5274), .CLK(clk), .Q(ram[837]) );
  DFFPOSX1 ram_reg_52__4_ ( .D(n5273), .CLK(clk), .Q(ram[836]) );
  DFFPOSX1 ram_reg_52__3_ ( .D(n5272), .CLK(clk), .Q(ram[835]) );
  DFFPOSX1 ram_reg_52__2_ ( .D(n5271), .CLK(clk), .Q(ram[834]) );
  DFFPOSX1 ram_reg_52__1_ ( .D(n5270), .CLK(clk), .Q(ram[833]) );
  DFFPOSX1 ram_reg_52__0_ ( .D(n5269), .CLK(clk), .Q(ram[832]) );
  DFFPOSX1 ram_reg_51__15_ ( .D(n5268), .CLK(clk), .Q(ram[831]) );
  DFFPOSX1 ram_reg_51__14_ ( .D(n5267), .CLK(clk), .Q(ram[830]) );
  DFFPOSX1 ram_reg_51__13_ ( .D(n5266), .CLK(clk), .Q(ram[829]) );
  DFFPOSX1 ram_reg_51__12_ ( .D(n5265), .CLK(clk), .Q(ram[828]) );
  DFFPOSX1 ram_reg_51__11_ ( .D(n5264), .CLK(clk), .Q(ram[827]) );
  DFFPOSX1 ram_reg_51__10_ ( .D(n5263), .CLK(clk), .Q(ram[826]) );
  DFFPOSX1 ram_reg_51__9_ ( .D(n5262), .CLK(clk), .Q(ram[825]) );
  DFFPOSX1 ram_reg_51__8_ ( .D(n5261), .CLK(clk), .Q(ram[824]) );
  DFFPOSX1 ram_reg_51__7_ ( .D(n5260), .CLK(clk), .Q(ram[823]) );
  DFFPOSX1 ram_reg_51__6_ ( .D(n5259), .CLK(clk), .Q(ram[822]) );
  DFFPOSX1 ram_reg_51__5_ ( .D(n5258), .CLK(clk), .Q(ram[821]) );
  DFFPOSX1 ram_reg_51__4_ ( .D(n5257), .CLK(clk), .Q(ram[820]) );
  DFFPOSX1 ram_reg_51__3_ ( .D(n5256), .CLK(clk), .Q(ram[819]) );
  DFFPOSX1 ram_reg_51__2_ ( .D(n5255), .CLK(clk), .Q(ram[818]) );
  DFFPOSX1 ram_reg_51__1_ ( .D(n5254), .CLK(clk), .Q(ram[817]) );
  DFFPOSX1 ram_reg_51__0_ ( .D(n5253), .CLK(clk), .Q(ram[816]) );
  DFFPOSX1 ram_reg_50__15_ ( .D(n5252), .CLK(clk), .Q(ram[815]) );
  DFFPOSX1 ram_reg_50__14_ ( .D(n5251), .CLK(clk), .Q(ram[814]) );
  DFFPOSX1 ram_reg_50__13_ ( .D(n5250), .CLK(clk), .Q(ram[813]) );
  DFFPOSX1 ram_reg_50__12_ ( .D(n5249), .CLK(clk), .Q(ram[812]) );
  DFFPOSX1 ram_reg_50__11_ ( .D(n5248), .CLK(clk), .Q(ram[811]) );
  DFFPOSX1 ram_reg_50__10_ ( .D(n5247), .CLK(clk), .Q(ram[810]) );
  DFFPOSX1 ram_reg_50__9_ ( .D(n5246), .CLK(clk), .Q(ram[809]) );
  DFFPOSX1 ram_reg_50__8_ ( .D(n5245), .CLK(clk), .Q(ram[808]) );
  DFFPOSX1 ram_reg_50__7_ ( .D(n5244), .CLK(clk), .Q(ram[807]) );
  DFFPOSX1 ram_reg_50__6_ ( .D(n5243), .CLK(clk), .Q(ram[806]) );
  DFFPOSX1 ram_reg_50__5_ ( .D(n5242), .CLK(clk), .Q(ram[805]) );
  DFFPOSX1 ram_reg_50__4_ ( .D(n5241), .CLK(clk), .Q(ram[804]) );
  DFFPOSX1 ram_reg_50__3_ ( .D(n5240), .CLK(clk), .Q(ram[803]) );
  DFFPOSX1 ram_reg_50__2_ ( .D(n5239), .CLK(clk), .Q(ram[802]) );
  DFFPOSX1 ram_reg_50__1_ ( .D(n5238), .CLK(clk), .Q(ram[801]) );
  DFFPOSX1 ram_reg_50__0_ ( .D(n5237), .CLK(clk), .Q(ram[800]) );
  DFFPOSX1 ram_reg_49__15_ ( .D(n5236), .CLK(clk), .Q(ram[799]) );
  DFFPOSX1 ram_reg_49__14_ ( .D(n5235), .CLK(clk), .Q(ram[798]) );
  DFFPOSX1 ram_reg_49__13_ ( .D(n5234), .CLK(clk), .Q(ram[797]) );
  DFFPOSX1 ram_reg_49__12_ ( .D(n5233), .CLK(clk), .Q(ram[796]) );
  DFFPOSX1 ram_reg_49__11_ ( .D(n5232), .CLK(clk), .Q(ram[795]) );
  DFFPOSX1 ram_reg_49__10_ ( .D(n5231), .CLK(clk), .Q(ram[794]) );
  DFFPOSX1 ram_reg_49__9_ ( .D(n5230), .CLK(clk), .Q(ram[793]) );
  DFFPOSX1 ram_reg_49__8_ ( .D(n5229), .CLK(clk), .Q(ram[792]) );
  DFFPOSX1 ram_reg_49__7_ ( .D(n5228), .CLK(clk), .Q(ram[791]) );
  DFFPOSX1 ram_reg_49__6_ ( .D(n5227), .CLK(clk), .Q(ram[790]) );
  DFFPOSX1 ram_reg_49__5_ ( .D(n5226), .CLK(clk), .Q(ram[789]) );
  DFFPOSX1 ram_reg_49__4_ ( .D(n5225), .CLK(clk), .Q(ram[788]) );
  DFFPOSX1 ram_reg_49__3_ ( .D(n5224), .CLK(clk), .Q(ram[787]) );
  DFFPOSX1 ram_reg_49__2_ ( .D(n5223), .CLK(clk), .Q(ram[786]) );
  DFFPOSX1 ram_reg_49__1_ ( .D(n5222), .CLK(clk), .Q(ram[785]) );
  DFFPOSX1 ram_reg_49__0_ ( .D(n5221), .CLK(clk), .Q(ram[784]) );
  DFFPOSX1 ram_reg_48__15_ ( .D(n5220), .CLK(clk), .Q(ram[783]) );
  DFFPOSX1 ram_reg_48__14_ ( .D(n5219), .CLK(clk), .Q(ram[782]) );
  DFFPOSX1 ram_reg_48__13_ ( .D(n5218), .CLK(clk), .Q(ram[781]) );
  DFFPOSX1 ram_reg_48__12_ ( .D(n5217), .CLK(clk), .Q(ram[780]) );
  DFFPOSX1 ram_reg_48__11_ ( .D(n5216), .CLK(clk), .Q(ram[779]) );
  DFFPOSX1 ram_reg_48__10_ ( .D(n5215), .CLK(clk), .Q(ram[778]) );
  DFFPOSX1 ram_reg_48__9_ ( .D(n5214), .CLK(clk), .Q(ram[777]) );
  DFFPOSX1 ram_reg_48__8_ ( .D(n5213), .CLK(clk), .Q(ram[776]) );
  DFFPOSX1 ram_reg_48__7_ ( .D(n5212), .CLK(clk), .Q(ram[775]) );
  DFFPOSX1 ram_reg_48__6_ ( .D(n5211), .CLK(clk), .Q(ram[774]) );
  DFFPOSX1 ram_reg_48__5_ ( .D(n5210), .CLK(clk), .Q(ram[773]) );
  DFFPOSX1 ram_reg_48__4_ ( .D(n5209), .CLK(clk), .Q(ram[772]) );
  DFFPOSX1 ram_reg_48__3_ ( .D(n5208), .CLK(clk), .Q(ram[771]) );
  DFFPOSX1 ram_reg_48__2_ ( .D(n5207), .CLK(clk), .Q(ram[770]) );
  DFFPOSX1 ram_reg_48__1_ ( .D(n5206), .CLK(clk), .Q(ram[769]) );
  DFFPOSX1 ram_reg_48__0_ ( .D(n5205), .CLK(clk), .Q(ram[768]) );
  DFFPOSX1 ram_reg_47__15_ ( .D(n5204), .CLK(clk), .Q(ram[767]) );
  DFFPOSX1 ram_reg_47__14_ ( .D(n5203), .CLK(clk), .Q(ram[766]) );
  DFFPOSX1 ram_reg_47__13_ ( .D(n5202), .CLK(clk), .Q(ram[765]) );
  DFFPOSX1 ram_reg_47__12_ ( .D(n5201), .CLK(clk), .Q(ram[764]) );
  DFFPOSX1 ram_reg_47__11_ ( .D(n5200), .CLK(clk), .Q(ram[763]) );
  DFFPOSX1 ram_reg_47__10_ ( .D(n5199), .CLK(clk), .Q(ram[762]) );
  DFFPOSX1 ram_reg_47__9_ ( .D(n5198), .CLK(clk), .Q(ram[761]) );
  DFFPOSX1 ram_reg_47__8_ ( .D(n5197), .CLK(clk), .Q(ram[760]) );
  DFFPOSX1 ram_reg_47__7_ ( .D(n5196), .CLK(clk), .Q(ram[759]) );
  DFFPOSX1 ram_reg_47__6_ ( .D(n5195), .CLK(clk), .Q(ram[758]) );
  DFFPOSX1 ram_reg_47__5_ ( .D(n5194), .CLK(clk), .Q(ram[757]) );
  DFFPOSX1 ram_reg_47__4_ ( .D(n5193), .CLK(clk), .Q(ram[756]) );
  DFFPOSX1 ram_reg_47__3_ ( .D(n5192), .CLK(clk), .Q(ram[755]) );
  DFFPOSX1 ram_reg_47__2_ ( .D(n5191), .CLK(clk), .Q(ram[754]) );
  DFFPOSX1 ram_reg_47__1_ ( .D(n5190), .CLK(clk), .Q(ram[753]) );
  DFFPOSX1 ram_reg_47__0_ ( .D(n5189), .CLK(clk), .Q(ram[752]) );
  DFFPOSX1 ram_reg_46__15_ ( .D(n5188), .CLK(clk), .Q(ram[751]) );
  DFFPOSX1 ram_reg_46__14_ ( .D(n5187), .CLK(clk), .Q(ram[750]) );
  DFFPOSX1 ram_reg_46__13_ ( .D(n5186), .CLK(clk), .Q(ram[749]) );
  DFFPOSX1 ram_reg_46__12_ ( .D(n5185), .CLK(clk), .Q(ram[748]) );
  DFFPOSX1 ram_reg_46__11_ ( .D(n5184), .CLK(clk), .Q(ram[747]) );
  DFFPOSX1 ram_reg_46__10_ ( .D(n5183), .CLK(clk), .Q(ram[746]) );
  DFFPOSX1 ram_reg_46__9_ ( .D(n5182), .CLK(clk), .Q(ram[745]) );
  DFFPOSX1 ram_reg_46__8_ ( .D(n5181), .CLK(clk), .Q(ram[744]) );
  DFFPOSX1 ram_reg_46__7_ ( .D(n5180), .CLK(clk), .Q(ram[743]) );
  DFFPOSX1 ram_reg_46__6_ ( .D(n5179), .CLK(clk), .Q(ram[742]) );
  DFFPOSX1 ram_reg_46__5_ ( .D(n5178), .CLK(clk), .Q(ram[741]) );
  DFFPOSX1 ram_reg_46__4_ ( .D(n5177), .CLK(clk), .Q(ram[740]) );
  DFFPOSX1 ram_reg_46__3_ ( .D(n5176), .CLK(clk), .Q(ram[739]) );
  DFFPOSX1 ram_reg_46__2_ ( .D(n5175), .CLK(clk), .Q(ram[738]) );
  DFFPOSX1 ram_reg_46__1_ ( .D(n5174), .CLK(clk), .Q(ram[737]) );
  DFFPOSX1 ram_reg_46__0_ ( .D(n5173), .CLK(clk), .Q(ram[736]) );
  DFFPOSX1 ram_reg_45__15_ ( .D(n5172), .CLK(clk), .Q(ram[735]) );
  DFFPOSX1 ram_reg_45__14_ ( .D(n5171), .CLK(clk), .Q(ram[734]) );
  DFFPOSX1 ram_reg_45__13_ ( .D(n5170), .CLK(clk), .Q(ram[733]) );
  DFFPOSX1 ram_reg_45__12_ ( .D(n5169), .CLK(clk), .Q(ram[732]) );
  DFFPOSX1 ram_reg_45__11_ ( .D(n5168), .CLK(clk), .Q(ram[731]) );
  DFFPOSX1 ram_reg_45__10_ ( .D(n5167), .CLK(clk), .Q(ram[730]) );
  DFFPOSX1 ram_reg_45__9_ ( .D(n5166), .CLK(clk), .Q(ram[729]) );
  DFFPOSX1 ram_reg_45__8_ ( .D(n5165), .CLK(clk), .Q(ram[728]) );
  DFFPOSX1 ram_reg_45__7_ ( .D(n5164), .CLK(clk), .Q(ram[727]) );
  DFFPOSX1 ram_reg_45__6_ ( .D(n5163), .CLK(clk), .Q(ram[726]) );
  DFFPOSX1 ram_reg_45__5_ ( .D(n5162), .CLK(clk), .Q(ram[725]) );
  DFFPOSX1 ram_reg_45__4_ ( .D(n5161), .CLK(clk), .Q(ram[724]) );
  DFFPOSX1 ram_reg_45__3_ ( .D(n5160), .CLK(clk), .Q(ram[723]) );
  DFFPOSX1 ram_reg_45__2_ ( .D(n5159), .CLK(clk), .Q(ram[722]) );
  DFFPOSX1 ram_reg_45__1_ ( .D(n5158), .CLK(clk), .Q(ram[721]) );
  DFFPOSX1 ram_reg_45__0_ ( .D(n5157), .CLK(clk), .Q(ram[720]) );
  DFFPOSX1 ram_reg_44__15_ ( .D(n5156), .CLK(clk), .Q(ram[719]) );
  DFFPOSX1 ram_reg_44__14_ ( .D(n5155), .CLK(clk), .Q(ram[718]) );
  DFFPOSX1 ram_reg_44__13_ ( .D(n5154), .CLK(clk), .Q(ram[717]) );
  DFFPOSX1 ram_reg_44__12_ ( .D(n5153), .CLK(clk), .Q(ram[716]) );
  DFFPOSX1 ram_reg_44__11_ ( .D(n5152), .CLK(clk), .Q(ram[715]) );
  DFFPOSX1 ram_reg_44__10_ ( .D(n5151), .CLK(clk), .Q(ram[714]) );
  DFFPOSX1 ram_reg_44__9_ ( .D(n5150), .CLK(clk), .Q(ram[713]) );
  DFFPOSX1 ram_reg_44__8_ ( .D(n5149), .CLK(clk), .Q(ram[712]) );
  DFFPOSX1 ram_reg_44__7_ ( .D(n5148), .CLK(clk), .Q(ram[711]) );
  DFFPOSX1 ram_reg_44__6_ ( .D(n5147), .CLK(clk), .Q(ram[710]) );
  DFFPOSX1 ram_reg_44__5_ ( .D(n5146), .CLK(clk), .Q(ram[709]) );
  DFFPOSX1 ram_reg_44__4_ ( .D(n5145), .CLK(clk), .Q(ram[708]) );
  DFFPOSX1 ram_reg_44__3_ ( .D(n5144), .CLK(clk), .Q(ram[707]) );
  DFFPOSX1 ram_reg_44__2_ ( .D(n5143), .CLK(clk), .Q(ram[706]) );
  DFFPOSX1 ram_reg_44__1_ ( .D(n5142), .CLK(clk), .Q(ram[705]) );
  DFFPOSX1 ram_reg_44__0_ ( .D(n5141), .CLK(clk), .Q(ram[704]) );
  DFFPOSX1 ram_reg_43__15_ ( .D(n5140), .CLK(clk), .Q(ram[703]) );
  DFFPOSX1 ram_reg_43__14_ ( .D(n5139), .CLK(clk), .Q(ram[702]) );
  DFFPOSX1 ram_reg_43__13_ ( .D(n5138), .CLK(clk), .Q(ram[701]) );
  DFFPOSX1 ram_reg_43__12_ ( .D(n5137), .CLK(clk), .Q(ram[700]) );
  DFFPOSX1 ram_reg_43__11_ ( .D(n5136), .CLK(clk), .Q(ram[699]) );
  DFFPOSX1 ram_reg_43__10_ ( .D(n5135), .CLK(clk), .Q(ram[698]) );
  DFFPOSX1 ram_reg_43__9_ ( .D(n5134), .CLK(clk), .Q(ram[697]) );
  DFFPOSX1 ram_reg_43__8_ ( .D(n5133), .CLK(clk), .Q(ram[696]) );
  DFFPOSX1 ram_reg_43__7_ ( .D(n5132), .CLK(clk), .Q(ram[695]) );
  DFFPOSX1 ram_reg_43__6_ ( .D(n5131), .CLK(clk), .Q(ram[694]) );
  DFFPOSX1 ram_reg_43__5_ ( .D(n5130), .CLK(clk), .Q(ram[693]) );
  DFFPOSX1 ram_reg_43__4_ ( .D(n5129), .CLK(clk), .Q(ram[692]) );
  DFFPOSX1 ram_reg_43__3_ ( .D(n5128), .CLK(clk), .Q(ram[691]) );
  DFFPOSX1 ram_reg_43__2_ ( .D(n5127), .CLK(clk), .Q(ram[690]) );
  DFFPOSX1 ram_reg_43__1_ ( .D(n5126), .CLK(clk), .Q(ram[689]) );
  DFFPOSX1 ram_reg_43__0_ ( .D(n5125), .CLK(clk), .Q(ram[688]) );
  DFFPOSX1 ram_reg_42__15_ ( .D(n5124), .CLK(clk), .Q(ram[687]) );
  DFFPOSX1 ram_reg_42__14_ ( .D(n5123), .CLK(clk), .Q(ram[686]) );
  DFFPOSX1 ram_reg_42__13_ ( .D(n5122), .CLK(clk), .Q(ram[685]) );
  DFFPOSX1 ram_reg_42__12_ ( .D(n5121), .CLK(clk), .Q(ram[684]) );
  DFFPOSX1 ram_reg_42__11_ ( .D(n5120), .CLK(clk), .Q(ram[683]) );
  DFFPOSX1 ram_reg_42__10_ ( .D(n5119), .CLK(clk), .Q(ram[682]) );
  DFFPOSX1 ram_reg_42__9_ ( .D(n5118), .CLK(clk), .Q(ram[681]) );
  DFFPOSX1 ram_reg_42__8_ ( .D(n5117), .CLK(clk), .Q(ram[680]) );
  DFFPOSX1 ram_reg_42__7_ ( .D(n5116), .CLK(clk), .Q(ram[679]) );
  DFFPOSX1 ram_reg_42__6_ ( .D(n5115), .CLK(clk), .Q(ram[678]) );
  DFFPOSX1 ram_reg_42__5_ ( .D(n5114), .CLK(clk), .Q(ram[677]) );
  DFFPOSX1 ram_reg_42__4_ ( .D(n5113), .CLK(clk), .Q(ram[676]) );
  DFFPOSX1 ram_reg_42__3_ ( .D(n5112), .CLK(clk), .Q(ram[675]) );
  DFFPOSX1 ram_reg_42__2_ ( .D(n5111), .CLK(clk), .Q(ram[674]) );
  DFFPOSX1 ram_reg_42__1_ ( .D(n5110), .CLK(clk), .Q(ram[673]) );
  DFFPOSX1 ram_reg_42__0_ ( .D(n5109), .CLK(clk), .Q(ram[672]) );
  DFFPOSX1 ram_reg_41__15_ ( .D(n5108), .CLK(clk), .Q(ram[671]) );
  DFFPOSX1 ram_reg_41__14_ ( .D(n5107), .CLK(clk), .Q(ram[670]) );
  DFFPOSX1 ram_reg_41__13_ ( .D(n5106), .CLK(clk), .Q(ram[669]) );
  DFFPOSX1 ram_reg_41__12_ ( .D(n5105), .CLK(clk), .Q(ram[668]) );
  DFFPOSX1 ram_reg_41__11_ ( .D(n5104), .CLK(clk), .Q(ram[667]) );
  DFFPOSX1 ram_reg_41__10_ ( .D(n5103), .CLK(clk), .Q(ram[666]) );
  DFFPOSX1 ram_reg_41__9_ ( .D(n5102), .CLK(clk), .Q(ram[665]) );
  DFFPOSX1 ram_reg_41__8_ ( .D(n5101), .CLK(clk), .Q(ram[664]) );
  DFFPOSX1 ram_reg_41__7_ ( .D(n5100), .CLK(clk), .Q(ram[663]) );
  DFFPOSX1 ram_reg_41__6_ ( .D(n5099), .CLK(clk), .Q(ram[662]) );
  DFFPOSX1 ram_reg_41__5_ ( .D(n5098), .CLK(clk), .Q(ram[661]) );
  DFFPOSX1 ram_reg_41__4_ ( .D(n5097), .CLK(clk), .Q(ram[660]) );
  DFFPOSX1 ram_reg_41__3_ ( .D(n5096), .CLK(clk), .Q(ram[659]) );
  DFFPOSX1 ram_reg_41__2_ ( .D(n5095), .CLK(clk), .Q(ram[658]) );
  DFFPOSX1 ram_reg_41__1_ ( .D(n5094), .CLK(clk), .Q(ram[657]) );
  DFFPOSX1 ram_reg_41__0_ ( .D(n5093), .CLK(clk), .Q(ram[656]) );
  DFFPOSX1 ram_reg_40__15_ ( .D(n5092), .CLK(clk), .Q(ram[655]) );
  DFFPOSX1 ram_reg_40__14_ ( .D(n5091), .CLK(clk), .Q(ram[654]) );
  DFFPOSX1 ram_reg_40__13_ ( .D(n5090), .CLK(clk), .Q(ram[653]) );
  DFFPOSX1 ram_reg_40__12_ ( .D(n5089), .CLK(clk), .Q(ram[652]) );
  DFFPOSX1 ram_reg_40__11_ ( .D(n5088), .CLK(clk), .Q(ram[651]) );
  DFFPOSX1 ram_reg_40__10_ ( .D(n5087), .CLK(clk), .Q(ram[650]) );
  DFFPOSX1 ram_reg_40__9_ ( .D(n5086), .CLK(clk), .Q(ram[649]) );
  DFFPOSX1 ram_reg_40__8_ ( .D(n5085), .CLK(clk), .Q(ram[648]) );
  DFFPOSX1 ram_reg_40__7_ ( .D(n5084), .CLK(clk), .Q(ram[647]) );
  DFFPOSX1 ram_reg_40__6_ ( .D(n5083), .CLK(clk), .Q(ram[646]) );
  DFFPOSX1 ram_reg_40__5_ ( .D(n5082), .CLK(clk), .Q(ram[645]) );
  DFFPOSX1 ram_reg_40__4_ ( .D(n5081), .CLK(clk), .Q(ram[644]) );
  DFFPOSX1 ram_reg_40__3_ ( .D(n5080), .CLK(clk), .Q(ram[643]) );
  DFFPOSX1 ram_reg_40__2_ ( .D(n5079), .CLK(clk), .Q(ram[642]) );
  DFFPOSX1 ram_reg_40__1_ ( .D(n5078), .CLK(clk), .Q(ram[641]) );
  DFFPOSX1 ram_reg_40__0_ ( .D(n5077), .CLK(clk), .Q(ram[640]) );
  DFFPOSX1 ram_reg_39__15_ ( .D(n5076), .CLK(clk), .Q(ram[639]) );
  DFFPOSX1 ram_reg_39__14_ ( .D(n5075), .CLK(clk), .Q(ram[638]) );
  DFFPOSX1 ram_reg_39__13_ ( .D(n5074), .CLK(clk), .Q(ram[637]) );
  DFFPOSX1 ram_reg_39__12_ ( .D(n5073), .CLK(clk), .Q(ram[636]) );
  DFFPOSX1 ram_reg_39__11_ ( .D(n5072), .CLK(clk), .Q(ram[635]) );
  DFFPOSX1 ram_reg_39__10_ ( .D(n5071), .CLK(clk), .Q(ram[634]) );
  DFFPOSX1 ram_reg_39__9_ ( .D(n5070), .CLK(clk), .Q(ram[633]) );
  DFFPOSX1 ram_reg_39__8_ ( .D(n5069), .CLK(clk), .Q(ram[632]) );
  DFFPOSX1 ram_reg_39__7_ ( .D(n5068), .CLK(clk), .Q(ram[631]) );
  DFFPOSX1 ram_reg_39__6_ ( .D(n5067), .CLK(clk), .Q(ram[630]) );
  DFFPOSX1 ram_reg_39__5_ ( .D(n5066), .CLK(clk), .Q(ram[629]) );
  DFFPOSX1 ram_reg_39__4_ ( .D(n5065), .CLK(clk), .Q(ram[628]) );
  DFFPOSX1 ram_reg_39__3_ ( .D(n5064), .CLK(clk), .Q(ram[627]) );
  DFFPOSX1 ram_reg_39__2_ ( .D(n5063), .CLK(clk), .Q(ram[626]) );
  DFFPOSX1 ram_reg_39__1_ ( .D(n5062), .CLK(clk), .Q(ram[625]) );
  DFFPOSX1 ram_reg_39__0_ ( .D(n5061), .CLK(clk), .Q(ram[624]) );
  DFFPOSX1 ram_reg_38__15_ ( .D(n5060), .CLK(clk), .Q(ram[623]) );
  DFFPOSX1 ram_reg_38__14_ ( .D(n5059), .CLK(clk), .Q(ram[622]) );
  DFFPOSX1 ram_reg_38__13_ ( .D(n5058), .CLK(clk), .Q(ram[621]) );
  DFFPOSX1 ram_reg_38__12_ ( .D(n5057), .CLK(clk), .Q(ram[620]) );
  DFFPOSX1 ram_reg_38__11_ ( .D(n5056), .CLK(clk), .Q(ram[619]) );
  DFFPOSX1 ram_reg_38__10_ ( .D(n5055), .CLK(clk), .Q(ram[618]) );
  DFFPOSX1 ram_reg_38__9_ ( .D(n5054), .CLK(clk), .Q(ram[617]) );
  DFFPOSX1 ram_reg_38__8_ ( .D(n5053), .CLK(clk), .Q(ram[616]) );
  DFFPOSX1 ram_reg_38__7_ ( .D(n5052), .CLK(clk), .Q(ram[615]) );
  DFFPOSX1 ram_reg_38__6_ ( .D(n5051), .CLK(clk), .Q(ram[614]) );
  DFFPOSX1 ram_reg_38__5_ ( .D(n5050), .CLK(clk), .Q(ram[613]) );
  DFFPOSX1 ram_reg_38__4_ ( .D(n5049), .CLK(clk), .Q(ram[612]) );
  DFFPOSX1 ram_reg_38__3_ ( .D(n5048), .CLK(clk), .Q(ram[611]) );
  DFFPOSX1 ram_reg_38__2_ ( .D(n5047), .CLK(clk), .Q(ram[610]) );
  DFFPOSX1 ram_reg_38__1_ ( .D(n5046), .CLK(clk), .Q(ram[609]) );
  DFFPOSX1 ram_reg_38__0_ ( .D(n5045), .CLK(clk), .Q(ram[608]) );
  DFFPOSX1 ram_reg_37__15_ ( .D(n5044), .CLK(clk), .Q(ram[607]) );
  DFFPOSX1 ram_reg_37__14_ ( .D(n5043), .CLK(clk), .Q(ram[606]) );
  DFFPOSX1 ram_reg_37__13_ ( .D(n5042), .CLK(clk), .Q(ram[605]) );
  DFFPOSX1 ram_reg_37__12_ ( .D(n5041), .CLK(clk), .Q(ram[604]) );
  DFFPOSX1 ram_reg_37__11_ ( .D(n5040), .CLK(clk), .Q(ram[603]) );
  DFFPOSX1 ram_reg_37__10_ ( .D(n5039), .CLK(clk), .Q(ram[602]) );
  DFFPOSX1 ram_reg_37__9_ ( .D(n5038), .CLK(clk), .Q(ram[601]) );
  DFFPOSX1 ram_reg_37__8_ ( .D(n5037), .CLK(clk), .Q(ram[600]) );
  DFFPOSX1 ram_reg_37__7_ ( .D(n5036), .CLK(clk), .Q(ram[599]) );
  DFFPOSX1 ram_reg_37__6_ ( .D(n5035), .CLK(clk), .Q(ram[598]) );
  DFFPOSX1 ram_reg_37__5_ ( .D(n5034), .CLK(clk), .Q(ram[597]) );
  DFFPOSX1 ram_reg_37__4_ ( .D(n5033), .CLK(clk), .Q(ram[596]) );
  DFFPOSX1 ram_reg_37__3_ ( .D(n5032), .CLK(clk), .Q(ram[595]) );
  DFFPOSX1 ram_reg_37__2_ ( .D(n5031), .CLK(clk), .Q(ram[594]) );
  DFFPOSX1 ram_reg_37__1_ ( .D(n5030), .CLK(clk), .Q(ram[593]) );
  DFFPOSX1 ram_reg_37__0_ ( .D(n5029), .CLK(clk), .Q(ram[592]) );
  DFFPOSX1 ram_reg_36__15_ ( .D(n5028), .CLK(clk), .Q(ram[591]) );
  DFFPOSX1 ram_reg_36__14_ ( .D(n5027), .CLK(clk), .Q(ram[590]) );
  DFFPOSX1 ram_reg_36__13_ ( .D(n5026), .CLK(clk), .Q(ram[589]) );
  DFFPOSX1 ram_reg_36__12_ ( .D(n5025), .CLK(clk), .Q(ram[588]) );
  DFFPOSX1 ram_reg_36__11_ ( .D(n5024), .CLK(clk), .Q(ram[587]) );
  DFFPOSX1 ram_reg_36__10_ ( .D(n5023), .CLK(clk), .Q(ram[586]) );
  DFFPOSX1 ram_reg_36__9_ ( .D(n5022), .CLK(clk), .Q(ram[585]) );
  DFFPOSX1 ram_reg_36__8_ ( .D(n5021), .CLK(clk), .Q(ram[584]) );
  DFFPOSX1 ram_reg_36__7_ ( .D(n5020), .CLK(clk), .Q(ram[583]) );
  DFFPOSX1 ram_reg_36__6_ ( .D(n5019), .CLK(clk), .Q(ram[582]) );
  DFFPOSX1 ram_reg_36__5_ ( .D(n5018), .CLK(clk), .Q(ram[581]) );
  DFFPOSX1 ram_reg_36__4_ ( .D(n5017), .CLK(clk), .Q(ram[580]) );
  DFFPOSX1 ram_reg_36__3_ ( .D(n5016), .CLK(clk), .Q(ram[579]) );
  DFFPOSX1 ram_reg_36__2_ ( .D(n5015), .CLK(clk), .Q(ram[578]) );
  DFFPOSX1 ram_reg_36__1_ ( .D(n5014), .CLK(clk), .Q(ram[577]) );
  DFFPOSX1 ram_reg_36__0_ ( .D(n5013), .CLK(clk), .Q(ram[576]) );
  DFFPOSX1 ram_reg_35__15_ ( .D(n5012), .CLK(clk), .Q(ram[575]) );
  DFFPOSX1 ram_reg_35__14_ ( .D(n5011), .CLK(clk), .Q(ram[574]) );
  DFFPOSX1 ram_reg_35__13_ ( .D(n5010), .CLK(clk), .Q(ram[573]) );
  DFFPOSX1 ram_reg_35__12_ ( .D(n5009), .CLK(clk), .Q(ram[572]) );
  DFFPOSX1 ram_reg_35__11_ ( .D(n5008), .CLK(clk), .Q(ram[571]) );
  DFFPOSX1 ram_reg_35__10_ ( .D(n5007), .CLK(clk), .Q(ram[570]) );
  DFFPOSX1 ram_reg_35__9_ ( .D(n5006), .CLK(clk), .Q(ram[569]) );
  DFFPOSX1 ram_reg_35__8_ ( .D(n5005), .CLK(clk), .Q(ram[568]) );
  DFFPOSX1 ram_reg_35__7_ ( .D(n5004), .CLK(clk), .Q(ram[567]) );
  DFFPOSX1 ram_reg_35__6_ ( .D(n5003), .CLK(clk), .Q(ram[566]) );
  DFFPOSX1 ram_reg_35__5_ ( .D(n5002), .CLK(clk), .Q(ram[565]) );
  DFFPOSX1 ram_reg_35__4_ ( .D(n5001), .CLK(clk), .Q(ram[564]) );
  DFFPOSX1 ram_reg_35__3_ ( .D(n5000), .CLK(clk), .Q(ram[563]) );
  DFFPOSX1 ram_reg_35__2_ ( .D(n4999), .CLK(clk), .Q(ram[562]) );
  DFFPOSX1 ram_reg_35__1_ ( .D(n4998), .CLK(clk), .Q(ram[561]) );
  DFFPOSX1 ram_reg_35__0_ ( .D(n4997), .CLK(clk), .Q(ram[560]) );
  DFFPOSX1 ram_reg_34__15_ ( .D(n4996), .CLK(clk), .Q(ram[559]) );
  DFFPOSX1 ram_reg_34__14_ ( .D(n4995), .CLK(clk), .Q(ram[558]) );
  DFFPOSX1 ram_reg_34__13_ ( .D(n4994), .CLK(clk), .Q(ram[557]) );
  DFFPOSX1 ram_reg_34__12_ ( .D(n4993), .CLK(clk), .Q(ram[556]) );
  DFFPOSX1 ram_reg_34__11_ ( .D(n4992), .CLK(clk), .Q(ram[555]) );
  DFFPOSX1 ram_reg_34__10_ ( .D(n4991), .CLK(clk), .Q(ram[554]) );
  DFFPOSX1 ram_reg_34__9_ ( .D(n4990), .CLK(clk), .Q(ram[553]) );
  DFFPOSX1 ram_reg_34__8_ ( .D(n4989), .CLK(clk), .Q(ram[552]) );
  DFFPOSX1 ram_reg_34__7_ ( .D(n4988), .CLK(clk), .Q(ram[551]) );
  DFFPOSX1 ram_reg_34__6_ ( .D(n4987), .CLK(clk), .Q(ram[550]) );
  DFFPOSX1 ram_reg_34__5_ ( .D(n4986), .CLK(clk), .Q(ram[549]) );
  DFFPOSX1 ram_reg_34__4_ ( .D(n4985), .CLK(clk), .Q(ram[548]) );
  DFFPOSX1 ram_reg_34__3_ ( .D(n4984), .CLK(clk), .Q(ram[547]) );
  DFFPOSX1 ram_reg_34__2_ ( .D(n4983), .CLK(clk), .Q(ram[546]) );
  DFFPOSX1 ram_reg_34__1_ ( .D(n4982), .CLK(clk), .Q(ram[545]) );
  DFFPOSX1 ram_reg_34__0_ ( .D(n4981), .CLK(clk), .Q(ram[544]) );
  DFFPOSX1 ram_reg_33__15_ ( .D(n4980), .CLK(clk), .Q(ram[543]) );
  DFFPOSX1 ram_reg_33__14_ ( .D(n4979), .CLK(clk), .Q(ram[542]) );
  DFFPOSX1 ram_reg_33__13_ ( .D(n4978), .CLK(clk), .Q(ram[541]) );
  DFFPOSX1 ram_reg_33__12_ ( .D(n4977), .CLK(clk), .Q(ram[540]) );
  DFFPOSX1 ram_reg_33__11_ ( .D(n4976), .CLK(clk), .Q(ram[539]) );
  DFFPOSX1 ram_reg_33__10_ ( .D(n4975), .CLK(clk), .Q(ram[538]) );
  DFFPOSX1 ram_reg_33__9_ ( .D(n4974), .CLK(clk), .Q(ram[537]) );
  DFFPOSX1 ram_reg_33__8_ ( .D(n4973), .CLK(clk), .Q(ram[536]) );
  DFFPOSX1 ram_reg_33__7_ ( .D(n4972), .CLK(clk), .Q(ram[535]) );
  DFFPOSX1 ram_reg_33__6_ ( .D(n4971), .CLK(clk), .Q(ram[534]) );
  DFFPOSX1 ram_reg_33__5_ ( .D(n4970), .CLK(clk), .Q(ram[533]) );
  DFFPOSX1 ram_reg_33__4_ ( .D(n4969), .CLK(clk), .Q(ram[532]) );
  DFFPOSX1 ram_reg_33__3_ ( .D(n4968), .CLK(clk), .Q(ram[531]) );
  DFFPOSX1 ram_reg_33__2_ ( .D(n4967), .CLK(clk), .Q(ram[530]) );
  DFFPOSX1 ram_reg_33__1_ ( .D(n4966), .CLK(clk), .Q(ram[529]) );
  DFFPOSX1 ram_reg_33__0_ ( .D(n4965), .CLK(clk), .Q(ram[528]) );
  DFFPOSX1 ram_reg_32__15_ ( .D(n4964), .CLK(clk), .Q(ram[527]) );
  DFFPOSX1 ram_reg_32__14_ ( .D(n4963), .CLK(clk), .Q(ram[526]) );
  DFFPOSX1 ram_reg_32__13_ ( .D(n4962), .CLK(clk), .Q(ram[525]) );
  DFFPOSX1 ram_reg_32__12_ ( .D(n4961), .CLK(clk), .Q(ram[524]) );
  DFFPOSX1 ram_reg_32__11_ ( .D(n4960), .CLK(clk), .Q(ram[523]) );
  DFFPOSX1 ram_reg_32__10_ ( .D(n4959), .CLK(clk), .Q(ram[522]) );
  DFFPOSX1 ram_reg_32__9_ ( .D(n4958), .CLK(clk), .Q(ram[521]) );
  DFFPOSX1 ram_reg_32__8_ ( .D(n4957), .CLK(clk), .Q(ram[520]) );
  DFFPOSX1 ram_reg_32__7_ ( .D(n4956), .CLK(clk), .Q(ram[519]) );
  DFFPOSX1 ram_reg_32__6_ ( .D(n4955), .CLK(clk), .Q(ram[518]) );
  DFFPOSX1 ram_reg_32__5_ ( .D(n4954), .CLK(clk), .Q(ram[517]) );
  DFFPOSX1 ram_reg_32__4_ ( .D(n4953), .CLK(clk), .Q(ram[516]) );
  DFFPOSX1 ram_reg_32__3_ ( .D(n4952), .CLK(clk), .Q(ram[515]) );
  DFFPOSX1 ram_reg_32__2_ ( .D(n4951), .CLK(clk), .Q(ram[514]) );
  DFFPOSX1 ram_reg_32__1_ ( .D(n4950), .CLK(clk), .Q(ram[513]) );
  DFFPOSX1 ram_reg_32__0_ ( .D(n4949), .CLK(clk), .Q(ram[512]) );
  DFFPOSX1 ram_reg_31__15_ ( .D(n4948), .CLK(clk), .Q(ram[511]) );
  DFFPOSX1 ram_reg_31__14_ ( .D(n4947), .CLK(clk), .Q(ram[510]) );
  DFFPOSX1 ram_reg_31__13_ ( .D(n4946), .CLK(clk), .Q(ram[509]) );
  DFFPOSX1 ram_reg_31__12_ ( .D(n4945), .CLK(clk), .Q(ram[508]) );
  DFFPOSX1 ram_reg_31__11_ ( .D(n4944), .CLK(clk), .Q(ram[507]) );
  DFFPOSX1 ram_reg_31__10_ ( .D(n4943), .CLK(clk), .Q(ram[506]) );
  DFFPOSX1 ram_reg_31__9_ ( .D(n4942), .CLK(clk), .Q(ram[505]) );
  DFFPOSX1 ram_reg_31__8_ ( .D(n4941), .CLK(clk), .Q(ram[504]) );
  DFFPOSX1 ram_reg_31__7_ ( .D(n4940), .CLK(clk), .Q(ram[503]) );
  DFFPOSX1 ram_reg_31__6_ ( .D(n4939), .CLK(clk), .Q(ram[502]) );
  DFFPOSX1 ram_reg_31__5_ ( .D(n4938), .CLK(clk), .Q(ram[501]) );
  DFFPOSX1 ram_reg_31__4_ ( .D(n4937), .CLK(clk), .Q(ram[500]) );
  DFFPOSX1 ram_reg_31__3_ ( .D(n4936), .CLK(clk), .Q(ram[499]) );
  DFFPOSX1 ram_reg_31__2_ ( .D(n4935), .CLK(clk), .Q(ram[498]) );
  DFFPOSX1 ram_reg_31__1_ ( .D(n4934), .CLK(clk), .Q(ram[497]) );
  DFFPOSX1 ram_reg_31__0_ ( .D(n4933), .CLK(clk), .Q(ram[496]) );
  DFFPOSX1 ram_reg_30__15_ ( .D(n4932), .CLK(clk), .Q(ram[495]) );
  DFFPOSX1 ram_reg_30__14_ ( .D(n4931), .CLK(clk), .Q(ram[494]) );
  DFFPOSX1 ram_reg_30__13_ ( .D(n4930), .CLK(clk), .Q(ram[493]) );
  DFFPOSX1 ram_reg_30__12_ ( .D(n4929), .CLK(clk), .Q(ram[492]) );
  DFFPOSX1 ram_reg_30__11_ ( .D(n4928), .CLK(clk), .Q(ram[491]) );
  DFFPOSX1 ram_reg_30__10_ ( .D(n4927), .CLK(clk), .Q(ram[490]) );
  DFFPOSX1 ram_reg_30__9_ ( .D(n4926), .CLK(clk), .Q(ram[489]) );
  DFFPOSX1 ram_reg_30__8_ ( .D(n4925), .CLK(clk), .Q(ram[488]) );
  DFFPOSX1 ram_reg_30__7_ ( .D(n4924), .CLK(clk), .Q(ram[487]) );
  DFFPOSX1 ram_reg_30__6_ ( .D(n4923), .CLK(clk), .Q(ram[486]) );
  DFFPOSX1 ram_reg_30__5_ ( .D(n4922), .CLK(clk), .Q(ram[485]) );
  DFFPOSX1 ram_reg_30__4_ ( .D(n4921), .CLK(clk), .Q(ram[484]) );
  DFFPOSX1 ram_reg_30__3_ ( .D(n4920), .CLK(clk), .Q(ram[483]) );
  DFFPOSX1 ram_reg_30__2_ ( .D(n4919), .CLK(clk), .Q(ram[482]) );
  DFFPOSX1 ram_reg_30__1_ ( .D(n4918), .CLK(clk), .Q(ram[481]) );
  DFFPOSX1 ram_reg_30__0_ ( .D(n4917), .CLK(clk), .Q(ram[480]) );
  DFFPOSX1 ram_reg_29__15_ ( .D(n4916), .CLK(clk), .Q(ram[479]) );
  DFFPOSX1 ram_reg_29__14_ ( .D(n4915), .CLK(clk), .Q(ram[478]) );
  DFFPOSX1 ram_reg_29__13_ ( .D(n4914), .CLK(clk), .Q(ram[477]) );
  DFFPOSX1 ram_reg_29__12_ ( .D(n4913), .CLK(clk), .Q(ram[476]) );
  DFFPOSX1 ram_reg_29__11_ ( .D(n4912), .CLK(clk), .Q(ram[475]) );
  DFFPOSX1 ram_reg_29__10_ ( .D(n4911), .CLK(clk), .Q(ram[474]) );
  DFFPOSX1 ram_reg_29__9_ ( .D(n4910), .CLK(clk), .Q(ram[473]) );
  DFFPOSX1 ram_reg_29__8_ ( .D(n4909), .CLK(clk), .Q(ram[472]) );
  DFFPOSX1 ram_reg_29__7_ ( .D(n4908), .CLK(clk), .Q(ram[471]) );
  DFFPOSX1 ram_reg_29__6_ ( .D(n4907), .CLK(clk), .Q(ram[470]) );
  DFFPOSX1 ram_reg_29__5_ ( .D(n4906), .CLK(clk), .Q(ram[469]) );
  DFFPOSX1 ram_reg_29__4_ ( .D(n4905), .CLK(clk), .Q(ram[468]) );
  DFFPOSX1 ram_reg_29__3_ ( .D(n4904), .CLK(clk), .Q(ram[467]) );
  DFFPOSX1 ram_reg_29__2_ ( .D(n4903), .CLK(clk), .Q(ram[466]) );
  DFFPOSX1 ram_reg_29__1_ ( .D(n4902), .CLK(clk), .Q(ram[465]) );
  DFFPOSX1 ram_reg_29__0_ ( .D(n4901), .CLK(clk), .Q(ram[464]) );
  DFFPOSX1 ram_reg_28__15_ ( .D(n4900), .CLK(clk), .Q(ram[463]) );
  DFFPOSX1 ram_reg_28__14_ ( .D(n4899), .CLK(clk), .Q(ram[462]) );
  DFFPOSX1 ram_reg_28__13_ ( .D(n4898), .CLK(clk), .Q(ram[461]) );
  DFFPOSX1 ram_reg_28__12_ ( .D(n4897), .CLK(clk), .Q(ram[460]) );
  DFFPOSX1 ram_reg_28__11_ ( .D(n4896), .CLK(clk), .Q(ram[459]) );
  DFFPOSX1 ram_reg_28__10_ ( .D(n4895), .CLK(clk), .Q(ram[458]) );
  DFFPOSX1 ram_reg_28__9_ ( .D(n4894), .CLK(clk), .Q(ram[457]) );
  DFFPOSX1 ram_reg_28__8_ ( .D(n4893), .CLK(clk), .Q(ram[456]) );
  DFFPOSX1 ram_reg_28__7_ ( .D(n4892), .CLK(clk), .Q(ram[455]) );
  DFFPOSX1 ram_reg_28__6_ ( .D(n4891), .CLK(clk), .Q(ram[454]) );
  DFFPOSX1 ram_reg_28__5_ ( .D(n4890), .CLK(clk), .Q(ram[453]) );
  DFFPOSX1 ram_reg_28__4_ ( .D(n4889), .CLK(clk), .Q(ram[452]) );
  DFFPOSX1 ram_reg_28__3_ ( .D(n4888), .CLK(clk), .Q(ram[451]) );
  DFFPOSX1 ram_reg_28__2_ ( .D(n4887), .CLK(clk), .Q(ram[450]) );
  DFFPOSX1 ram_reg_28__1_ ( .D(n4886), .CLK(clk), .Q(ram[449]) );
  DFFPOSX1 ram_reg_28__0_ ( .D(n4885), .CLK(clk), .Q(ram[448]) );
  DFFPOSX1 ram_reg_27__15_ ( .D(n4884), .CLK(clk), .Q(ram[447]) );
  DFFPOSX1 ram_reg_27__14_ ( .D(n4883), .CLK(clk), .Q(ram[446]) );
  DFFPOSX1 ram_reg_27__13_ ( .D(n4882), .CLK(clk), .Q(ram[445]) );
  DFFPOSX1 ram_reg_27__12_ ( .D(n4881), .CLK(clk), .Q(ram[444]) );
  DFFPOSX1 ram_reg_27__11_ ( .D(n4880), .CLK(clk), .Q(ram[443]) );
  DFFPOSX1 ram_reg_27__10_ ( .D(n4879), .CLK(clk), .Q(ram[442]) );
  DFFPOSX1 ram_reg_27__9_ ( .D(n4878), .CLK(clk), .Q(ram[441]) );
  DFFPOSX1 ram_reg_27__8_ ( .D(n4877), .CLK(clk), .Q(ram[440]) );
  DFFPOSX1 ram_reg_27__7_ ( .D(n4876), .CLK(clk), .Q(ram[439]) );
  DFFPOSX1 ram_reg_27__6_ ( .D(n4875), .CLK(clk), .Q(ram[438]) );
  DFFPOSX1 ram_reg_27__5_ ( .D(n4874), .CLK(clk), .Q(ram[437]) );
  DFFPOSX1 ram_reg_27__4_ ( .D(n4873), .CLK(clk), .Q(ram[436]) );
  DFFPOSX1 ram_reg_27__3_ ( .D(n4872), .CLK(clk), .Q(ram[435]) );
  DFFPOSX1 ram_reg_27__2_ ( .D(n4871), .CLK(clk), .Q(ram[434]) );
  DFFPOSX1 ram_reg_27__1_ ( .D(n4870), .CLK(clk), .Q(ram[433]) );
  DFFPOSX1 ram_reg_27__0_ ( .D(n4869), .CLK(clk), .Q(ram[432]) );
  DFFPOSX1 ram_reg_26__15_ ( .D(n4868), .CLK(clk), .Q(ram[431]) );
  DFFPOSX1 ram_reg_26__14_ ( .D(n4867), .CLK(clk), .Q(ram[430]) );
  DFFPOSX1 ram_reg_26__13_ ( .D(n4866), .CLK(clk), .Q(ram[429]) );
  DFFPOSX1 ram_reg_26__12_ ( .D(n4865), .CLK(clk), .Q(ram[428]) );
  DFFPOSX1 ram_reg_26__11_ ( .D(n4864), .CLK(clk), .Q(ram[427]) );
  DFFPOSX1 ram_reg_26__10_ ( .D(n4863), .CLK(clk), .Q(ram[426]) );
  DFFPOSX1 ram_reg_26__9_ ( .D(n4862), .CLK(clk), .Q(ram[425]) );
  DFFPOSX1 ram_reg_26__8_ ( .D(n4861), .CLK(clk), .Q(ram[424]) );
  DFFPOSX1 ram_reg_26__7_ ( .D(n4860), .CLK(clk), .Q(ram[423]) );
  DFFPOSX1 ram_reg_26__6_ ( .D(n4859), .CLK(clk), .Q(ram[422]) );
  DFFPOSX1 ram_reg_26__5_ ( .D(n4858), .CLK(clk), .Q(ram[421]) );
  DFFPOSX1 ram_reg_26__4_ ( .D(n4857), .CLK(clk), .Q(ram[420]) );
  DFFPOSX1 ram_reg_26__3_ ( .D(n4856), .CLK(clk), .Q(ram[419]) );
  DFFPOSX1 ram_reg_26__2_ ( .D(n4855), .CLK(clk), .Q(ram[418]) );
  DFFPOSX1 ram_reg_26__1_ ( .D(n4854), .CLK(clk), .Q(ram[417]) );
  DFFPOSX1 ram_reg_26__0_ ( .D(n4853), .CLK(clk), .Q(ram[416]) );
  DFFPOSX1 ram_reg_25__15_ ( .D(n4852), .CLK(clk), .Q(ram[415]) );
  DFFPOSX1 ram_reg_25__14_ ( .D(n4851), .CLK(clk), .Q(ram[414]) );
  DFFPOSX1 ram_reg_25__13_ ( .D(n4850), .CLK(clk), .Q(ram[413]) );
  DFFPOSX1 ram_reg_25__12_ ( .D(n4849), .CLK(clk), .Q(ram[412]) );
  DFFPOSX1 ram_reg_25__11_ ( .D(n4848), .CLK(clk), .Q(ram[411]) );
  DFFPOSX1 ram_reg_25__10_ ( .D(n4847), .CLK(clk), .Q(ram[410]) );
  DFFPOSX1 ram_reg_25__9_ ( .D(n4846), .CLK(clk), .Q(ram[409]) );
  DFFPOSX1 ram_reg_25__8_ ( .D(n4845), .CLK(clk), .Q(ram[408]) );
  DFFPOSX1 ram_reg_25__7_ ( .D(n4844), .CLK(clk), .Q(ram[407]) );
  DFFPOSX1 ram_reg_25__6_ ( .D(n4843), .CLK(clk), .Q(ram[406]) );
  DFFPOSX1 ram_reg_25__5_ ( .D(n4842), .CLK(clk), .Q(ram[405]) );
  DFFPOSX1 ram_reg_25__4_ ( .D(n4841), .CLK(clk), .Q(ram[404]) );
  DFFPOSX1 ram_reg_25__3_ ( .D(n4840), .CLK(clk), .Q(ram[403]) );
  DFFPOSX1 ram_reg_25__2_ ( .D(n4839), .CLK(clk), .Q(ram[402]) );
  DFFPOSX1 ram_reg_25__1_ ( .D(n4838), .CLK(clk), .Q(ram[401]) );
  DFFPOSX1 ram_reg_25__0_ ( .D(n4837), .CLK(clk), .Q(ram[400]) );
  DFFPOSX1 ram_reg_24__15_ ( .D(n4836), .CLK(clk), .Q(ram[399]) );
  DFFPOSX1 ram_reg_24__14_ ( .D(n4835), .CLK(clk), .Q(ram[398]) );
  DFFPOSX1 ram_reg_24__13_ ( .D(n4834), .CLK(clk), .Q(ram[397]) );
  DFFPOSX1 ram_reg_24__12_ ( .D(n4833), .CLK(clk), .Q(ram[396]) );
  DFFPOSX1 ram_reg_24__11_ ( .D(n4832), .CLK(clk), .Q(ram[395]) );
  DFFPOSX1 ram_reg_24__10_ ( .D(n4831), .CLK(clk), .Q(ram[394]) );
  DFFPOSX1 ram_reg_24__9_ ( .D(n4830), .CLK(clk), .Q(ram[393]) );
  DFFPOSX1 ram_reg_24__8_ ( .D(n4829), .CLK(clk), .Q(ram[392]) );
  DFFPOSX1 ram_reg_24__7_ ( .D(n4828), .CLK(clk), .Q(ram[391]) );
  DFFPOSX1 ram_reg_24__6_ ( .D(n4827), .CLK(clk), .Q(ram[390]) );
  DFFPOSX1 ram_reg_24__5_ ( .D(n4826), .CLK(clk), .Q(ram[389]) );
  DFFPOSX1 ram_reg_24__4_ ( .D(n4825), .CLK(clk), .Q(ram[388]) );
  DFFPOSX1 ram_reg_24__3_ ( .D(n4824), .CLK(clk), .Q(ram[387]) );
  DFFPOSX1 ram_reg_24__2_ ( .D(n4823), .CLK(clk), .Q(ram[386]) );
  DFFPOSX1 ram_reg_24__1_ ( .D(n4822), .CLK(clk), .Q(ram[385]) );
  DFFPOSX1 ram_reg_24__0_ ( .D(n4821), .CLK(clk), .Q(ram[384]) );
  DFFPOSX1 ram_reg_23__15_ ( .D(n4820), .CLK(clk), .Q(ram[383]) );
  DFFPOSX1 ram_reg_23__14_ ( .D(n4819), .CLK(clk), .Q(ram[382]) );
  DFFPOSX1 ram_reg_23__13_ ( .D(n4818), .CLK(clk), .Q(ram[381]) );
  DFFPOSX1 ram_reg_23__12_ ( .D(n4817), .CLK(clk), .Q(ram[380]) );
  DFFPOSX1 ram_reg_23__11_ ( .D(n4816), .CLK(clk), .Q(ram[379]) );
  DFFPOSX1 ram_reg_23__10_ ( .D(n4815), .CLK(clk), .Q(ram[378]) );
  DFFPOSX1 ram_reg_23__9_ ( .D(n4814), .CLK(clk), .Q(ram[377]) );
  DFFPOSX1 ram_reg_23__8_ ( .D(n4813), .CLK(clk), .Q(ram[376]) );
  DFFPOSX1 ram_reg_23__7_ ( .D(n4812), .CLK(clk), .Q(ram[375]) );
  DFFPOSX1 ram_reg_23__6_ ( .D(n4811), .CLK(clk), .Q(ram[374]) );
  DFFPOSX1 ram_reg_23__5_ ( .D(n4810), .CLK(clk), .Q(ram[373]) );
  DFFPOSX1 ram_reg_23__4_ ( .D(n4809), .CLK(clk), .Q(ram[372]) );
  DFFPOSX1 ram_reg_23__3_ ( .D(n4808), .CLK(clk), .Q(ram[371]) );
  DFFPOSX1 ram_reg_23__2_ ( .D(n4807), .CLK(clk), .Q(ram[370]) );
  DFFPOSX1 ram_reg_23__1_ ( .D(n4806), .CLK(clk), .Q(ram[369]) );
  DFFPOSX1 ram_reg_23__0_ ( .D(n4805), .CLK(clk), .Q(ram[368]) );
  DFFPOSX1 ram_reg_22__15_ ( .D(n4804), .CLK(clk), .Q(ram[367]) );
  DFFPOSX1 ram_reg_22__14_ ( .D(n4803), .CLK(clk), .Q(ram[366]) );
  DFFPOSX1 ram_reg_22__13_ ( .D(n4802), .CLK(clk), .Q(ram[365]) );
  DFFPOSX1 ram_reg_22__12_ ( .D(n4801), .CLK(clk), .Q(ram[364]) );
  DFFPOSX1 ram_reg_22__11_ ( .D(n4800), .CLK(clk), .Q(ram[363]) );
  DFFPOSX1 ram_reg_22__10_ ( .D(n4799), .CLK(clk), .Q(ram[362]) );
  DFFPOSX1 ram_reg_22__9_ ( .D(n4798), .CLK(clk), .Q(ram[361]) );
  DFFPOSX1 ram_reg_22__8_ ( .D(n4797), .CLK(clk), .Q(ram[360]) );
  DFFPOSX1 ram_reg_22__7_ ( .D(n4796), .CLK(clk), .Q(ram[359]) );
  DFFPOSX1 ram_reg_22__6_ ( .D(n4795), .CLK(clk), .Q(ram[358]) );
  DFFPOSX1 ram_reg_22__5_ ( .D(n4794), .CLK(clk), .Q(ram[357]) );
  DFFPOSX1 ram_reg_22__4_ ( .D(n4793), .CLK(clk), .Q(ram[356]) );
  DFFPOSX1 ram_reg_22__3_ ( .D(n4792), .CLK(clk), .Q(ram[355]) );
  DFFPOSX1 ram_reg_22__2_ ( .D(n4791), .CLK(clk), .Q(ram[354]) );
  DFFPOSX1 ram_reg_22__1_ ( .D(n4790), .CLK(clk), .Q(ram[353]) );
  DFFPOSX1 ram_reg_22__0_ ( .D(n4789), .CLK(clk), .Q(ram[352]) );
  DFFPOSX1 ram_reg_21__15_ ( .D(n4788), .CLK(clk), .Q(ram[351]) );
  DFFPOSX1 ram_reg_21__14_ ( .D(n4787), .CLK(clk), .Q(ram[350]) );
  DFFPOSX1 ram_reg_21__13_ ( .D(n4786), .CLK(clk), .Q(ram[349]) );
  DFFPOSX1 ram_reg_21__12_ ( .D(n4785), .CLK(clk), .Q(ram[348]) );
  DFFPOSX1 ram_reg_21__11_ ( .D(n4784), .CLK(clk), .Q(ram[347]) );
  DFFPOSX1 ram_reg_21__10_ ( .D(n4783), .CLK(clk), .Q(ram[346]) );
  DFFPOSX1 ram_reg_21__9_ ( .D(n4782), .CLK(clk), .Q(ram[345]) );
  DFFPOSX1 ram_reg_21__8_ ( .D(n4781), .CLK(clk), .Q(ram[344]) );
  DFFPOSX1 ram_reg_21__7_ ( .D(n4780), .CLK(clk), .Q(ram[343]) );
  DFFPOSX1 ram_reg_21__6_ ( .D(n4779), .CLK(clk), .Q(ram[342]) );
  DFFPOSX1 ram_reg_21__5_ ( .D(n4778), .CLK(clk), .Q(ram[341]) );
  DFFPOSX1 ram_reg_21__4_ ( .D(n4777), .CLK(clk), .Q(ram[340]) );
  DFFPOSX1 ram_reg_21__3_ ( .D(n4776), .CLK(clk), .Q(ram[339]) );
  DFFPOSX1 ram_reg_21__2_ ( .D(n4775), .CLK(clk), .Q(ram[338]) );
  DFFPOSX1 ram_reg_21__1_ ( .D(n4774), .CLK(clk), .Q(ram[337]) );
  DFFPOSX1 ram_reg_21__0_ ( .D(n4773), .CLK(clk), .Q(ram[336]) );
  DFFPOSX1 ram_reg_20__15_ ( .D(n4772), .CLK(clk), .Q(ram[335]) );
  DFFPOSX1 ram_reg_20__14_ ( .D(n4771), .CLK(clk), .Q(ram[334]) );
  DFFPOSX1 ram_reg_20__13_ ( .D(n4770), .CLK(clk), .Q(ram[333]) );
  DFFPOSX1 ram_reg_20__12_ ( .D(n4769), .CLK(clk), .Q(ram[332]) );
  DFFPOSX1 ram_reg_20__11_ ( .D(n4768), .CLK(clk), .Q(ram[331]) );
  DFFPOSX1 ram_reg_20__10_ ( .D(n4767), .CLK(clk), .Q(ram[330]) );
  DFFPOSX1 ram_reg_20__9_ ( .D(n4766), .CLK(clk), .Q(ram[329]) );
  DFFPOSX1 ram_reg_20__8_ ( .D(n4765), .CLK(clk), .Q(ram[328]) );
  DFFPOSX1 ram_reg_20__7_ ( .D(n4764), .CLK(clk), .Q(ram[327]) );
  DFFPOSX1 ram_reg_20__6_ ( .D(n4763), .CLK(clk), .Q(ram[326]) );
  DFFPOSX1 ram_reg_20__5_ ( .D(n4762), .CLK(clk), .Q(ram[325]) );
  DFFPOSX1 ram_reg_20__4_ ( .D(n4761), .CLK(clk), .Q(ram[324]) );
  DFFPOSX1 ram_reg_20__3_ ( .D(n4760), .CLK(clk), .Q(ram[323]) );
  DFFPOSX1 ram_reg_20__2_ ( .D(n4759), .CLK(clk), .Q(ram[322]) );
  DFFPOSX1 ram_reg_20__1_ ( .D(n4758), .CLK(clk), .Q(ram[321]) );
  DFFPOSX1 ram_reg_20__0_ ( .D(n4757), .CLK(clk), .Q(ram[320]) );
  DFFPOSX1 ram_reg_19__15_ ( .D(n4756), .CLK(clk), .Q(ram[319]) );
  DFFPOSX1 ram_reg_19__14_ ( .D(n4755), .CLK(clk), .Q(ram[318]) );
  DFFPOSX1 ram_reg_19__13_ ( .D(n4754), .CLK(clk), .Q(ram[317]) );
  DFFPOSX1 ram_reg_19__12_ ( .D(n4753), .CLK(clk), .Q(ram[316]) );
  DFFPOSX1 ram_reg_19__11_ ( .D(n4752), .CLK(clk), .Q(ram[315]) );
  DFFPOSX1 ram_reg_19__10_ ( .D(n4751), .CLK(clk), .Q(ram[314]) );
  DFFPOSX1 ram_reg_19__9_ ( .D(n4750), .CLK(clk), .Q(ram[313]) );
  DFFPOSX1 ram_reg_19__8_ ( .D(n4749), .CLK(clk), .Q(ram[312]) );
  DFFPOSX1 ram_reg_19__7_ ( .D(n4748), .CLK(clk), .Q(ram[311]) );
  DFFPOSX1 ram_reg_19__6_ ( .D(n4747), .CLK(clk), .Q(ram[310]) );
  DFFPOSX1 ram_reg_19__5_ ( .D(n4746), .CLK(clk), .Q(ram[309]) );
  DFFPOSX1 ram_reg_19__4_ ( .D(n4745), .CLK(clk), .Q(ram[308]) );
  DFFPOSX1 ram_reg_19__3_ ( .D(n4744), .CLK(clk), .Q(ram[307]) );
  DFFPOSX1 ram_reg_19__2_ ( .D(n4743), .CLK(clk), .Q(ram[306]) );
  DFFPOSX1 ram_reg_19__1_ ( .D(n4742), .CLK(clk), .Q(ram[305]) );
  DFFPOSX1 ram_reg_19__0_ ( .D(n4741), .CLK(clk), .Q(ram[304]) );
  DFFPOSX1 ram_reg_18__15_ ( .D(n4740), .CLK(clk), .Q(ram[303]) );
  DFFPOSX1 ram_reg_18__14_ ( .D(n4739), .CLK(clk), .Q(ram[302]) );
  DFFPOSX1 ram_reg_18__13_ ( .D(n4738), .CLK(clk), .Q(ram[301]) );
  DFFPOSX1 ram_reg_18__12_ ( .D(n4737), .CLK(clk), .Q(ram[300]) );
  DFFPOSX1 ram_reg_18__11_ ( .D(n4736), .CLK(clk), .Q(ram[299]) );
  DFFPOSX1 ram_reg_18__10_ ( .D(n4735), .CLK(clk), .Q(ram[298]) );
  DFFPOSX1 ram_reg_18__9_ ( .D(n4734), .CLK(clk), .Q(ram[297]) );
  DFFPOSX1 ram_reg_18__8_ ( .D(n4733), .CLK(clk), .Q(ram[296]) );
  DFFPOSX1 ram_reg_18__7_ ( .D(n4732), .CLK(clk), .Q(ram[295]) );
  DFFPOSX1 ram_reg_18__6_ ( .D(n4731), .CLK(clk), .Q(ram[294]) );
  DFFPOSX1 ram_reg_18__5_ ( .D(n4730), .CLK(clk), .Q(ram[293]) );
  DFFPOSX1 ram_reg_18__4_ ( .D(n4729), .CLK(clk), .Q(ram[292]) );
  DFFPOSX1 ram_reg_18__3_ ( .D(n4728), .CLK(clk), .Q(ram[291]) );
  DFFPOSX1 ram_reg_18__2_ ( .D(n4727), .CLK(clk), .Q(ram[290]) );
  DFFPOSX1 ram_reg_18__1_ ( .D(n4726), .CLK(clk), .Q(ram[289]) );
  DFFPOSX1 ram_reg_18__0_ ( .D(n4725), .CLK(clk), .Q(ram[288]) );
  DFFPOSX1 ram_reg_17__15_ ( .D(n4724), .CLK(clk), .Q(ram[287]) );
  DFFPOSX1 ram_reg_17__14_ ( .D(n4723), .CLK(clk), .Q(ram[286]) );
  DFFPOSX1 ram_reg_17__13_ ( .D(n4722), .CLK(clk), .Q(ram[285]) );
  DFFPOSX1 ram_reg_17__12_ ( .D(n4721), .CLK(clk), .Q(ram[284]) );
  DFFPOSX1 ram_reg_17__11_ ( .D(n4720), .CLK(clk), .Q(ram[283]) );
  DFFPOSX1 ram_reg_17__10_ ( .D(n4719), .CLK(clk), .Q(ram[282]) );
  DFFPOSX1 ram_reg_17__9_ ( .D(n4718), .CLK(clk), .Q(ram[281]) );
  DFFPOSX1 ram_reg_17__8_ ( .D(n4717), .CLK(clk), .Q(ram[280]) );
  DFFPOSX1 ram_reg_17__7_ ( .D(n4716), .CLK(clk), .Q(ram[279]) );
  DFFPOSX1 ram_reg_17__6_ ( .D(n4715), .CLK(clk), .Q(ram[278]) );
  DFFPOSX1 ram_reg_17__5_ ( .D(n4714), .CLK(clk), .Q(ram[277]) );
  DFFPOSX1 ram_reg_17__4_ ( .D(n4713), .CLK(clk), .Q(ram[276]) );
  DFFPOSX1 ram_reg_17__3_ ( .D(n4712), .CLK(clk), .Q(ram[275]) );
  DFFPOSX1 ram_reg_17__2_ ( .D(n4711), .CLK(clk), .Q(ram[274]) );
  DFFPOSX1 ram_reg_17__1_ ( .D(n4710), .CLK(clk), .Q(ram[273]) );
  DFFPOSX1 ram_reg_17__0_ ( .D(n4709), .CLK(clk), .Q(ram[272]) );
  DFFPOSX1 ram_reg_16__15_ ( .D(n4708), .CLK(clk), .Q(ram[271]) );
  DFFPOSX1 ram_reg_16__14_ ( .D(n4707), .CLK(clk), .Q(ram[270]) );
  DFFPOSX1 ram_reg_16__13_ ( .D(n4706), .CLK(clk), .Q(ram[269]) );
  DFFPOSX1 ram_reg_16__12_ ( .D(n4705), .CLK(clk), .Q(ram[268]) );
  DFFPOSX1 ram_reg_16__11_ ( .D(n4704), .CLK(clk), .Q(ram[267]) );
  DFFPOSX1 ram_reg_16__10_ ( .D(n4703), .CLK(clk), .Q(ram[266]) );
  DFFPOSX1 ram_reg_16__9_ ( .D(n4702), .CLK(clk), .Q(ram[265]) );
  DFFPOSX1 ram_reg_16__8_ ( .D(n4701), .CLK(clk), .Q(ram[264]) );
  DFFPOSX1 ram_reg_16__7_ ( .D(n4700), .CLK(clk), .Q(ram[263]) );
  DFFPOSX1 ram_reg_16__6_ ( .D(n4699), .CLK(clk), .Q(ram[262]) );
  DFFPOSX1 ram_reg_16__5_ ( .D(n4698), .CLK(clk), .Q(ram[261]) );
  DFFPOSX1 ram_reg_16__4_ ( .D(n4697), .CLK(clk), .Q(ram[260]) );
  DFFPOSX1 ram_reg_16__3_ ( .D(n4696), .CLK(clk), .Q(ram[259]) );
  DFFPOSX1 ram_reg_16__2_ ( .D(n4695), .CLK(clk), .Q(ram[258]) );
  DFFPOSX1 ram_reg_16__1_ ( .D(n4694), .CLK(clk), .Q(ram[257]) );
  DFFPOSX1 ram_reg_16__0_ ( .D(n4693), .CLK(clk), .Q(ram[256]) );
  DFFPOSX1 ram_reg_15__15_ ( .D(n4692), .CLK(clk), .Q(ram[255]) );
  DFFPOSX1 ram_reg_15__14_ ( .D(n4691), .CLK(clk), .Q(ram[254]) );
  DFFPOSX1 ram_reg_15__13_ ( .D(n4690), .CLK(clk), .Q(ram[253]) );
  DFFPOSX1 ram_reg_15__12_ ( .D(n4689), .CLK(clk), .Q(ram[252]) );
  DFFPOSX1 ram_reg_15__11_ ( .D(n4688), .CLK(clk), .Q(ram[251]) );
  DFFPOSX1 ram_reg_15__10_ ( .D(n4687), .CLK(clk), .Q(ram[250]) );
  DFFPOSX1 ram_reg_15__9_ ( .D(n4686), .CLK(clk), .Q(ram[249]) );
  DFFPOSX1 ram_reg_15__8_ ( .D(n4685), .CLK(clk), .Q(ram[248]) );
  DFFPOSX1 ram_reg_15__7_ ( .D(n4684), .CLK(clk), .Q(ram[247]) );
  DFFPOSX1 ram_reg_15__6_ ( .D(n4683), .CLK(clk), .Q(ram[246]) );
  DFFPOSX1 ram_reg_15__5_ ( .D(n4682), .CLK(clk), .Q(ram[245]) );
  DFFPOSX1 ram_reg_15__4_ ( .D(n4681), .CLK(clk), .Q(ram[244]) );
  DFFPOSX1 ram_reg_15__3_ ( .D(n4680), .CLK(clk), .Q(ram[243]) );
  DFFPOSX1 ram_reg_15__2_ ( .D(n4679), .CLK(clk), .Q(ram[242]) );
  DFFPOSX1 ram_reg_15__1_ ( .D(n4678), .CLK(clk), .Q(ram[241]) );
  DFFPOSX1 ram_reg_15__0_ ( .D(n4677), .CLK(clk), .Q(ram[240]) );
  DFFPOSX1 ram_reg_14__15_ ( .D(n4676), .CLK(clk), .Q(ram[239]) );
  DFFPOSX1 ram_reg_14__14_ ( .D(n4675), .CLK(clk), .Q(ram[238]) );
  DFFPOSX1 ram_reg_14__13_ ( .D(n4674), .CLK(clk), .Q(ram[237]) );
  DFFPOSX1 ram_reg_14__12_ ( .D(n4673), .CLK(clk), .Q(ram[236]) );
  DFFPOSX1 ram_reg_14__11_ ( .D(n4672), .CLK(clk), .Q(ram[235]) );
  DFFPOSX1 ram_reg_14__10_ ( .D(n4671), .CLK(clk), .Q(ram[234]) );
  DFFPOSX1 ram_reg_14__9_ ( .D(n4670), .CLK(clk), .Q(ram[233]) );
  DFFPOSX1 ram_reg_14__8_ ( .D(n4669), .CLK(clk), .Q(ram[232]) );
  DFFPOSX1 ram_reg_14__7_ ( .D(n4668), .CLK(clk), .Q(ram[231]) );
  DFFPOSX1 ram_reg_14__6_ ( .D(n4667), .CLK(clk), .Q(ram[230]) );
  DFFPOSX1 ram_reg_14__5_ ( .D(n4666), .CLK(clk), .Q(ram[229]) );
  DFFPOSX1 ram_reg_14__4_ ( .D(n4665), .CLK(clk), .Q(ram[228]) );
  DFFPOSX1 ram_reg_14__3_ ( .D(n4664), .CLK(clk), .Q(ram[227]) );
  DFFPOSX1 ram_reg_14__2_ ( .D(n4663), .CLK(clk), .Q(ram[226]) );
  DFFPOSX1 ram_reg_14__1_ ( .D(n4662), .CLK(clk), .Q(ram[225]) );
  DFFPOSX1 ram_reg_14__0_ ( .D(n4661), .CLK(clk), .Q(ram[224]) );
  DFFPOSX1 ram_reg_13__15_ ( .D(n4660), .CLK(clk), .Q(ram[223]) );
  DFFPOSX1 ram_reg_13__14_ ( .D(n4659), .CLK(clk), .Q(ram[222]) );
  DFFPOSX1 ram_reg_13__13_ ( .D(n4658), .CLK(clk), .Q(ram[221]) );
  DFFPOSX1 ram_reg_13__12_ ( .D(n4657), .CLK(clk), .Q(ram[220]) );
  DFFPOSX1 ram_reg_13__11_ ( .D(n4656), .CLK(clk), .Q(ram[219]) );
  DFFPOSX1 ram_reg_13__10_ ( .D(n4655), .CLK(clk), .Q(ram[218]) );
  DFFPOSX1 ram_reg_13__9_ ( .D(n4654), .CLK(clk), .Q(ram[217]) );
  DFFPOSX1 ram_reg_13__8_ ( .D(n4653), .CLK(clk), .Q(ram[216]) );
  DFFPOSX1 ram_reg_13__7_ ( .D(n4652), .CLK(clk), .Q(ram[215]) );
  DFFPOSX1 ram_reg_13__6_ ( .D(n4651), .CLK(clk), .Q(ram[214]) );
  DFFPOSX1 ram_reg_13__5_ ( .D(n4650), .CLK(clk), .Q(ram[213]) );
  DFFPOSX1 ram_reg_13__4_ ( .D(n4649), .CLK(clk), .Q(ram[212]) );
  DFFPOSX1 ram_reg_13__3_ ( .D(n4648), .CLK(clk), .Q(ram[211]) );
  DFFPOSX1 ram_reg_13__2_ ( .D(n4647), .CLK(clk), .Q(ram[210]) );
  DFFPOSX1 ram_reg_13__1_ ( .D(n4646), .CLK(clk), .Q(ram[209]) );
  DFFPOSX1 ram_reg_13__0_ ( .D(n4645), .CLK(clk), .Q(ram[208]) );
  DFFPOSX1 ram_reg_12__15_ ( .D(n4644), .CLK(clk), .Q(ram[207]) );
  DFFPOSX1 ram_reg_12__14_ ( .D(n4643), .CLK(clk), .Q(ram[206]) );
  DFFPOSX1 ram_reg_12__13_ ( .D(n4642), .CLK(clk), .Q(ram[205]) );
  DFFPOSX1 ram_reg_12__12_ ( .D(n4641), .CLK(clk), .Q(ram[204]) );
  DFFPOSX1 ram_reg_12__11_ ( .D(n4640), .CLK(clk), .Q(ram[203]) );
  DFFPOSX1 ram_reg_12__10_ ( .D(n4639), .CLK(clk), .Q(ram[202]) );
  DFFPOSX1 ram_reg_12__9_ ( .D(n4638), .CLK(clk), .Q(ram[201]) );
  DFFPOSX1 ram_reg_12__8_ ( .D(n4637), .CLK(clk), .Q(ram[200]) );
  DFFPOSX1 ram_reg_12__7_ ( .D(n4636), .CLK(clk), .Q(ram[199]) );
  DFFPOSX1 ram_reg_12__6_ ( .D(n4635), .CLK(clk), .Q(ram[198]) );
  DFFPOSX1 ram_reg_12__5_ ( .D(n4634), .CLK(clk), .Q(ram[197]) );
  DFFPOSX1 ram_reg_12__4_ ( .D(n4633), .CLK(clk), .Q(ram[196]) );
  DFFPOSX1 ram_reg_12__3_ ( .D(n4632), .CLK(clk), .Q(ram[195]) );
  DFFPOSX1 ram_reg_12__2_ ( .D(n4631), .CLK(clk), .Q(ram[194]) );
  DFFPOSX1 ram_reg_12__1_ ( .D(n4630), .CLK(clk), .Q(ram[193]) );
  DFFPOSX1 ram_reg_12__0_ ( .D(n4629), .CLK(clk), .Q(ram[192]) );
  DFFPOSX1 ram_reg_11__15_ ( .D(n4628), .CLK(clk), .Q(ram[191]) );
  DFFPOSX1 ram_reg_11__14_ ( .D(n4627), .CLK(clk), .Q(ram[190]) );
  DFFPOSX1 ram_reg_11__13_ ( .D(n4626), .CLK(clk), .Q(ram[189]) );
  DFFPOSX1 ram_reg_11__12_ ( .D(n4625), .CLK(clk), .Q(ram[188]) );
  DFFPOSX1 ram_reg_11__11_ ( .D(n4624), .CLK(clk), .Q(ram[187]) );
  DFFPOSX1 ram_reg_11__10_ ( .D(n4623), .CLK(clk), .Q(ram[186]) );
  DFFPOSX1 ram_reg_11__9_ ( .D(n4622), .CLK(clk), .Q(ram[185]) );
  DFFPOSX1 ram_reg_11__8_ ( .D(n4621), .CLK(clk), .Q(ram[184]) );
  DFFPOSX1 ram_reg_11__7_ ( .D(n4620), .CLK(clk), .Q(ram[183]) );
  DFFPOSX1 ram_reg_11__6_ ( .D(n4619), .CLK(clk), .Q(ram[182]) );
  DFFPOSX1 ram_reg_11__5_ ( .D(n4618), .CLK(clk), .Q(ram[181]) );
  DFFPOSX1 ram_reg_11__4_ ( .D(n4617), .CLK(clk), .Q(ram[180]) );
  DFFPOSX1 ram_reg_11__3_ ( .D(n4616), .CLK(clk), .Q(ram[179]) );
  DFFPOSX1 ram_reg_11__2_ ( .D(n4615), .CLK(clk), .Q(ram[178]) );
  DFFPOSX1 ram_reg_11__1_ ( .D(n4614), .CLK(clk), .Q(ram[177]) );
  DFFPOSX1 ram_reg_11__0_ ( .D(n4613), .CLK(clk), .Q(ram[176]) );
  DFFPOSX1 ram_reg_10__15_ ( .D(n4612), .CLK(clk), .Q(ram[175]) );
  DFFPOSX1 ram_reg_10__14_ ( .D(n4611), .CLK(clk), .Q(ram[174]) );
  DFFPOSX1 ram_reg_10__13_ ( .D(n4610), .CLK(clk), .Q(ram[173]) );
  DFFPOSX1 ram_reg_10__12_ ( .D(n4609), .CLK(clk), .Q(ram[172]) );
  DFFPOSX1 ram_reg_10__11_ ( .D(n4608), .CLK(clk), .Q(ram[171]) );
  DFFPOSX1 ram_reg_10__10_ ( .D(n4607), .CLK(clk), .Q(ram[170]) );
  DFFPOSX1 ram_reg_10__9_ ( .D(n4606), .CLK(clk), .Q(ram[169]) );
  DFFPOSX1 ram_reg_10__8_ ( .D(n4605), .CLK(clk), .Q(ram[168]) );
  DFFPOSX1 ram_reg_10__7_ ( .D(n4604), .CLK(clk), .Q(ram[167]) );
  DFFPOSX1 ram_reg_10__6_ ( .D(n4603), .CLK(clk), .Q(ram[166]) );
  DFFPOSX1 ram_reg_10__5_ ( .D(n4602), .CLK(clk), .Q(ram[165]) );
  DFFPOSX1 ram_reg_10__4_ ( .D(n4601), .CLK(clk), .Q(ram[164]) );
  DFFPOSX1 ram_reg_10__3_ ( .D(n4600), .CLK(clk), .Q(ram[163]) );
  DFFPOSX1 ram_reg_10__2_ ( .D(n4599), .CLK(clk), .Q(ram[162]) );
  DFFPOSX1 ram_reg_10__1_ ( .D(n4598), .CLK(clk), .Q(ram[161]) );
  DFFPOSX1 ram_reg_10__0_ ( .D(n4597), .CLK(clk), .Q(ram[160]) );
  DFFPOSX1 ram_reg_9__15_ ( .D(n4596), .CLK(clk), .Q(ram[159]) );
  DFFPOSX1 ram_reg_9__14_ ( .D(n4595), .CLK(clk), .Q(ram[158]) );
  DFFPOSX1 ram_reg_9__13_ ( .D(n4594), .CLK(clk), .Q(ram[157]) );
  DFFPOSX1 ram_reg_9__12_ ( .D(n4593), .CLK(clk), .Q(ram[156]) );
  DFFPOSX1 ram_reg_9__11_ ( .D(n4592), .CLK(clk), .Q(ram[155]) );
  DFFPOSX1 ram_reg_9__10_ ( .D(n4591), .CLK(clk), .Q(ram[154]) );
  DFFPOSX1 ram_reg_9__9_ ( .D(n4590), .CLK(clk), .Q(ram[153]) );
  DFFPOSX1 ram_reg_9__8_ ( .D(n4589), .CLK(clk), .Q(ram[152]) );
  DFFPOSX1 ram_reg_9__7_ ( .D(n4588), .CLK(clk), .Q(ram[151]) );
  DFFPOSX1 ram_reg_9__6_ ( .D(n4587), .CLK(clk), .Q(ram[150]) );
  DFFPOSX1 ram_reg_9__5_ ( .D(n4586), .CLK(clk), .Q(ram[149]) );
  DFFPOSX1 ram_reg_9__4_ ( .D(n4585), .CLK(clk), .Q(ram[148]) );
  DFFPOSX1 ram_reg_9__3_ ( .D(n4584), .CLK(clk), .Q(ram[147]) );
  DFFPOSX1 ram_reg_9__2_ ( .D(n4583), .CLK(clk), .Q(ram[146]) );
  DFFPOSX1 ram_reg_9__1_ ( .D(n4582), .CLK(clk), .Q(ram[145]) );
  DFFPOSX1 ram_reg_9__0_ ( .D(n4581), .CLK(clk), .Q(ram[144]) );
  DFFPOSX1 ram_reg_8__15_ ( .D(n4580), .CLK(clk), .Q(ram[143]) );
  DFFPOSX1 ram_reg_8__14_ ( .D(n4579), .CLK(clk), .Q(ram[142]) );
  DFFPOSX1 ram_reg_8__13_ ( .D(n4578), .CLK(clk), .Q(ram[141]) );
  DFFPOSX1 ram_reg_8__12_ ( .D(n4577), .CLK(clk), .Q(ram[140]) );
  DFFPOSX1 ram_reg_8__11_ ( .D(n4576), .CLK(clk), .Q(ram[139]) );
  DFFPOSX1 ram_reg_8__10_ ( .D(n4575), .CLK(clk), .Q(ram[138]) );
  DFFPOSX1 ram_reg_8__9_ ( .D(n4574), .CLK(clk), .Q(ram[137]) );
  DFFPOSX1 ram_reg_8__8_ ( .D(n4573), .CLK(clk), .Q(ram[136]) );
  DFFPOSX1 ram_reg_8__7_ ( .D(n4572), .CLK(clk), .Q(ram[135]) );
  DFFPOSX1 ram_reg_8__6_ ( .D(n4571), .CLK(clk), .Q(ram[134]) );
  DFFPOSX1 ram_reg_8__5_ ( .D(n4570), .CLK(clk), .Q(ram[133]) );
  DFFPOSX1 ram_reg_8__4_ ( .D(n4569), .CLK(clk), .Q(ram[132]) );
  DFFPOSX1 ram_reg_8__3_ ( .D(n4568), .CLK(clk), .Q(ram[131]) );
  DFFPOSX1 ram_reg_8__2_ ( .D(n4567), .CLK(clk), .Q(ram[130]) );
  DFFPOSX1 ram_reg_8__1_ ( .D(n4566), .CLK(clk), .Q(ram[129]) );
  DFFPOSX1 ram_reg_8__0_ ( .D(n4565), .CLK(clk), .Q(ram[128]) );
  DFFPOSX1 ram_reg_7__15_ ( .D(n4564), .CLK(clk), .Q(ram[127]) );
  DFFPOSX1 ram_reg_7__14_ ( .D(n4563), .CLK(clk), .Q(ram[126]) );
  DFFPOSX1 ram_reg_7__13_ ( .D(n4562), .CLK(clk), .Q(ram[125]) );
  DFFPOSX1 ram_reg_7__12_ ( .D(n4561), .CLK(clk), .Q(ram[124]) );
  DFFPOSX1 ram_reg_7__11_ ( .D(n4560), .CLK(clk), .Q(ram[123]) );
  DFFPOSX1 ram_reg_7__10_ ( .D(n4559), .CLK(clk), .Q(ram[122]) );
  DFFPOSX1 ram_reg_7__9_ ( .D(n4558), .CLK(clk), .Q(ram[121]) );
  DFFPOSX1 ram_reg_7__8_ ( .D(n4557), .CLK(clk), .Q(ram[120]) );
  DFFPOSX1 ram_reg_7__7_ ( .D(n4556), .CLK(clk), .Q(ram[119]) );
  DFFPOSX1 ram_reg_7__6_ ( .D(n4555), .CLK(clk), .Q(ram[118]) );
  DFFPOSX1 ram_reg_7__5_ ( .D(n4554), .CLK(clk), .Q(ram[117]) );
  DFFPOSX1 ram_reg_7__4_ ( .D(n4553), .CLK(clk), .Q(ram[116]) );
  DFFPOSX1 ram_reg_7__3_ ( .D(n4552), .CLK(clk), .Q(ram[115]) );
  DFFPOSX1 ram_reg_7__2_ ( .D(n4551), .CLK(clk), .Q(ram[114]) );
  DFFPOSX1 ram_reg_7__1_ ( .D(n4550), .CLK(clk), .Q(ram[113]) );
  DFFPOSX1 ram_reg_7__0_ ( .D(n4549), .CLK(clk), .Q(ram[112]) );
  DFFPOSX1 ram_reg_6__15_ ( .D(n4548), .CLK(clk), .Q(ram[111]) );
  DFFPOSX1 ram_reg_6__14_ ( .D(n4547), .CLK(clk), .Q(ram[110]) );
  DFFPOSX1 ram_reg_6__13_ ( .D(n4546), .CLK(clk), .Q(ram[109]) );
  DFFPOSX1 ram_reg_6__12_ ( .D(n4545), .CLK(clk), .Q(ram[108]) );
  DFFPOSX1 ram_reg_6__11_ ( .D(n4544), .CLK(clk), .Q(ram[107]) );
  DFFPOSX1 ram_reg_6__10_ ( .D(n4543), .CLK(clk), .Q(ram[106]) );
  DFFPOSX1 ram_reg_6__9_ ( .D(n4542), .CLK(clk), .Q(ram[105]) );
  DFFPOSX1 ram_reg_6__8_ ( .D(n4541), .CLK(clk), .Q(ram[104]) );
  DFFPOSX1 ram_reg_6__7_ ( .D(n4540), .CLK(clk), .Q(ram[103]) );
  DFFPOSX1 ram_reg_6__6_ ( .D(n4539), .CLK(clk), .Q(ram[102]) );
  DFFPOSX1 ram_reg_6__5_ ( .D(n4538), .CLK(clk), .Q(ram[101]) );
  DFFPOSX1 ram_reg_6__4_ ( .D(n4537), .CLK(clk), .Q(ram[100]) );
  DFFPOSX1 ram_reg_6__3_ ( .D(n4536), .CLK(clk), .Q(ram[99]) );
  DFFPOSX1 ram_reg_6__2_ ( .D(n4535), .CLK(clk), .Q(ram[98]) );
  DFFPOSX1 ram_reg_6__1_ ( .D(n4534), .CLK(clk), .Q(ram[97]) );
  DFFPOSX1 ram_reg_6__0_ ( .D(n4533), .CLK(clk), .Q(ram[96]) );
  DFFPOSX1 ram_reg_5__15_ ( .D(n4532), .CLK(clk), .Q(ram[95]) );
  DFFPOSX1 ram_reg_5__14_ ( .D(n4531), .CLK(clk), .Q(ram[94]) );
  DFFPOSX1 ram_reg_5__13_ ( .D(n4530), .CLK(clk), .Q(ram[93]) );
  DFFPOSX1 ram_reg_5__12_ ( .D(n4529), .CLK(clk), .Q(ram[92]) );
  DFFPOSX1 ram_reg_5__11_ ( .D(n4528), .CLK(clk), .Q(ram[91]) );
  DFFPOSX1 ram_reg_5__10_ ( .D(n4527), .CLK(clk), .Q(ram[90]) );
  DFFPOSX1 ram_reg_5__9_ ( .D(n4526), .CLK(clk), .Q(ram[89]) );
  DFFPOSX1 ram_reg_5__8_ ( .D(n4525), .CLK(clk), .Q(ram[88]) );
  DFFPOSX1 ram_reg_5__7_ ( .D(n4524), .CLK(clk), .Q(ram[87]) );
  DFFPOSX1 ram_reg_5__6_ ( .D(n4523), .CLK(clk), .Q(ram[86]) );
  DFFPOSX1 ram_reg_5__5_ ( .D(n4522), .CLK(clk), .Q(ram[85]) );
  DFFPOSX1 ram_reg_5__4_ ( .D(n4521), .CLK(clk), .Q(ram[84]) );
  DFFPOSX1 ram_reg_5__3_ ( .D(n4520), .CLK(clk), .Q(ram[83]) );
  DFFPOSX1 ram_reg_5__2_ ( .D(n4519), .CLK(clk), .Q(ram[82]) );
  DFFPOSX1 ram_reg_5__1_ ( .D(n4518), .CLK(clk), .Q(ram[81]) );
  DFFPOSX1 ram_reg_5__0_ ( .D(n4517), .CLK(clk), .Q(ram[80]) );
  DFFPOSX1 ram_reg_4__15_ ( .D(n4516), .CLK(clk), .Q(ram[79]) );
  DFFPOSX1 ram_reg_4__14_ ( .D(n4515), .CLK(clk), .Q(ram[78]) );
  DFFPOSX1 ram_reg_4__13_ ( .D(n4514), .CLK(clk), .Q(ram[77]) );
  DFFPOSX1 ram_reg_4__12_ ( .D(n4513), .CLK(clk), .Q(ram[76]) );
  DFFPOSX1 ram_reg_4__11_ ( .D(n4512), .CLK(clk), .Q(ram[75]) );
  DFFPOSX1 ram_reg_4__10_ ( .D(n4511), .CLK(clk), .Q(ram[74]) );
  DFFPOSX1 ram_reg_4__9_ ( .D(n4510), .CLK(clk), .Q(ram[73]) );
  DFFPOSX1 ram_reg_4__8_ ( .D(n4509), .CLK(clk), .Q(ram[72]) );
  DFFPOSX1 ram_reg_4__7_ ( .D(n4508), .CLK(clk), .Q(ram[71]) );
  DFFPOSX1 ram_reg_4__6_ ( .D(n4507), .CLK(clk), .Q(ram[70]) );
  DFFPOSX1 ram_reg_4__5_ ( .D(n4506), .CLK(clk), .Q(ram[69]) );
  DFFPOSX1 ram_reg_4__4_ ( .D(n4505), .CLK(clk), .Q(ram[68]) );
  DFFPOSX1 ram_reg_4__3_ ( .D(n4504), .CLK(clk), .Q(ram[67]) );
  DFFPOSX1 ram_reg_4__2_ ( .D(n4503), .CLK(clk), .Q(ram[66]) );
  DFFPOSX1 ram_reg_4__1_ ( .D(n4502), .CLK(clk), .Q(ram[65]) );
  DFFPOSX1 ram_reg_4__0_ ( .D(n4501), .CLK(clk), .Q(ram[64]) );
  DFFPOSX1 ram_reg_3__15_ ( .D(n4500), .CLK(clk), .Q(ram[63]) );
  DFFPOSX1 ram_reg_3__14_ ( .D(n4499), .CLK(clk), .Q(ram[62]) );
  DFFPOSX1 ram_reg_3__13_ ( .D(n4498), .CLK(clk), .Q(ram[61]) );
  DFFPOSX1 ram_reg_3__12_ ( .D(n4497), .CLK(clk), .Q(ram[60]) );
  DFFPOSX1 ram_reg_3__11_ ( .D(n4496), .CLK(clk), .Q(ram[59]) );
  DFFPOSX1 ram_reg_3__10_ ( .D(n4495), .CLK(clk), .Q(ram[58]) );
  DFFPOSX1 ram_reg_3__9_ ( .D(n4494), .CLK(clk), .Q(ram[57]) );
  DFFPOSX1 ram_reg_3__8_ ( .D(n4493), .CLK(clk), .Q(ram[56]) );
  DFFPOSX1 ram_reg_3__7_ ( .D(n4492), .CLK(clk), .Q(ram[55]) );
  DFFPOSX1 ram_reg_3__6_ ( .D(n4491), .CLK(clk), .Q(ram[54]) );
  DFFPOSX1 ram_reg_3__5_ ( .D(n4490), .CLK(clk), .Q(ram[53]) );
  DFFPOSX1 ram_reg_3__4_ ( .D(n4489), .CLK(clk), .Q(ram[52]) );
  DFFPOSX1 ram_reg_3__3_ ( .D(n4488), .CLK(clk), .Q(ram[51]) );
  DFFPOSX1 ram_reg_3__2_ ( .D(n4487), .CLK(clk), .Q(ram[50]) );
  DFFPOSX1 ram_reg_3__1_ ( .D(n4486), .CLK(clk), .Q(ram[49]) );
  DFFPOSX1 ram_reg_3__0_ ( .D(n4485), .CLK(clk), .Q(ram[48]) );
  DFFPOSX1 ram_reg_2__15_ ( .D(n4484), .CLK(clk), .Q(ram[47]) );
  DFFPOSX1 ram_reg_2__14_ ( .D(n4483), .CLK(clk), .Q(ram[46]) );
  DFFPOSX1 ram_reg_2__13_ ( .D(n4482), .CLK(clk), .Q(ram[45]) );
  DFFPOSX1 ram_reg_2__12_ ( .D(n4481), .CLK(clk), .Q(ram[44]) );
  DFFPOSX1 ram_reg_2__11_ ( .D(n4480), .CLK(clk), .Q(ram[43]) );
  DFFPOSX1 ram_reg_2__10_ ( .D(n4479), .CLK(clk), .Q(ram[42]) );
  DFFPOSX1 ram_reg_2__9_ ( .D(n4478), .CLK(clk), .Q(ram[41]) );
  DFFPOSX1 ram_reg_2__8_ ( .D(n4477), .CLK(clk), .Q(ram[40]) );
  DFFPOSX1 ram_reg_2__7_ ( .D(n4476), .CLK(clk), .Q(ram[39]) );
  DFFPOSX1 ram_reg_2__6_ ( .D(n4475), .CLK(clk), .Q(ram[38]) );
  DFFPOSX1 ram_reg_2__5_ ( .D(n4474), .CLK(clk), .Q(ram[37]) );
  DFFPOSX1 ram_reg_2__4_ ( .D(n4473), .CLK(clk), .Q(ram[36]) );
  DFFPOSX1 ram_reg_2__3_ ( .D(n4472), .CLK(clk), .Q(ram[35]) );
  DFFPOSX1 ram_reg_2__2_ ( .D(n4471), .CLK(clk), .Q(ram[34]) );
  DFFPOSX1 ram_reg_2__1_ ( .D(n4470), .CLK(clk), .Q(ram[33]) );
  DFFPOSX1 ram_reg_2__0_ ( .D(n4469), .CLK(clk), .Q(ram[32]) );
  DFFPOSX1 ram_reg_1__15_ ( .D(n4468), .CLK(clk), .Q(ram[31]) );
  DFFPOSX1 ram_reg_1__14_ ( .D(n4467), .CLK(clk), .Q(ram[30]) );
  DFFPOSX1 ram_reg_1__13_ ( .D(n4466), .CLK(clk), .Q(ram[29]) );
  DFFPOSX1 ram_reg_1__12_ ( .D(n4465), .CLK(clk), .Q(ram[28]) );
  DFFPOSX1 ram_reg_1__11_ ( .D(n4464), .CLK(clk), .Q(ram[27]) );
  DFFPOSX1 ram_reg_1__10_ ( .D(n4463), .CLK(clk), .Q(ram[26]) );
  DFFPOSX1 ram_reg_1__9_ ( .D(n4462), .CLK(clk), .Q(ram[25]) );
  DFFPOSX1 ram_reg_1__8_ ( .D(n4461), .CLK(clk), .Q(ram[24]) );
  DFFPOSX1 ram_reg_1__7_ ( .D(n4460), .CLK(clk), .Q(ram[23]) );
  DFFPOSX1 ram_reg_1__6_ ( .D(n4459), .CLK(clk), .Q(ram[22]) );
  DFFPOSX1 ram_reg_1__5_ ( .D(n4458), .CLK(clk), .Q(ram[21]) );
  DFFPOSX1 ram_reg_1__4_ ( .D(n4457), .CLK(clk), .Q(ram[20]) );
  DFFPOSX1 ram_reg_1__3_ ( .D(n4456), .CLK(clk), .Q(ram[19]) );
  DFFPOSX1 ram_reg_1__2_ ( .D(n4455), .CLK(clk), .Q(ram[18]) );
  DFFPOSX1 ram_reg_1__1_ ( .D(n4454), .CLK(clk), .Q(ram[17]) );
  DFFPOSX1 ram_reg_1__0_ ( .D(n4453), .CLK(clk), .Q(ram[16]) );
  DFFPOSX1 ram_reg_0__15_ ( .D(n4452), .CLK(clk), .Q(ram[15]) );
  DFFPOSX1 ram_reg_0__14_ ( .D(n4451), .CLK(clk), .Q(ram[14]) );
  DFFPOSX1 ram_reg_0__13_ ( .D(n4450), .CLK(clk), .Q(ram[13]) );
  DFFPOSX1 ram_reg_0__12_ ( .D(n4449), .CLK(clk), .Q(ram[12]) );
  DFFPOSX1 ram_reg_0__11_ ( .D(n4448), .CLK(clk), .Q(ram[11]) );
  DFFPOSX1 ram_reg_0__10_ ( .D(n4447), .CLK(clk), .Q(ram[10]) );
  DFFPOSX1 ram_reg_0__9_ ( .D(n4446), .CLK(clk), .Q(ram[9]) );
  DFFPOSX1 ram_reg_0__8_ ( .D(n4445), .CLK(clk), .Q(ram[8]) );
  DFFPOSX1 ram_reg_0__7_ ( .D(n4444), .CLK(clk), .Q(ram[7]) );
  DFFPOSX1 ram_reg_0__6_ ( .D(n4443), .CLK(clk), .Q(ram[6]) );
  DFFPOSX1 ram_reg_0__5_ ( .D(n4442), .CLK(clk), .Q(ram[5]) );
  DFFPOSX1 ram_reg_0__4_ ( .D(n4441), .CLK(clk), .Q(ram[4]) );
  DFFPOSX1 ram_reg_0__3_ ( .D(n4440), .CLK(clk), .Q(ram[3]) );
  DFFPOSX1 ram_reg_0__2_ ( .D(n4439), .CLK(clk), .Q(ram[2]) );
  DFFPOSX1 ram_reg_0__1_ ( .D(n4438), .CLK(clk), .Q(ram[1]) );
  DFFPOSX1 ram_reg_0__0_ ( .D(n4437), .CLK(clk), .Q(ram[0]) );
  OAI21X1 U38 ( .A(n13035), .B(n12776), .C(n38), .Y(n4437) );
  NAND2X1 U39 ( .A(ram[0]), .B(n13035), .Y(n38) );
  OAI21X1 U40 ( .A(n13035), .B(n12770), .C(n39), .Y(n4438) );
  NAND2X1 U41 ( .A(ram[1]), .B(n13035), .Y(n39) );
  OAI21X1 U42 ( .A(n13035), .B(n12762), .C(n40), .Y(n4439) );
  NAND2X1 U43 ( .A(ram[2]), .B(n13035), .Y(n40) );
  OAI21X1 U44 ( .A(n13035), .B(n12756), .C(n41), .Y(n4440) );
  NAND2X1 U45 ( .A(ram[3]), .B(n13035), .Y(n41) );
  OAI21X1 U46 ( .A(n13035), .B(n12750), .C(n42), .Y(n4441) );
  NAND2X1 U47 ( .A(ram[4]), .B(n13035), .Y(n42) );
  OAI21X1 U48 ( .A(n13035), .B(n12744), .C(n43), .Y(n4442) );
  NAND2X1 U49 ( .A(ram[5]), .B(n13035), .Y(n43) );
  OAI21X1 U50 ( .A(n13035), .B(n12738), .C(n44), .Y(n4443) );
  NAND2X1 U51 ( .A(ram[6]), .B(n13035), .Y(n44) );
  OAI21X1 U52 ( .A(n13035), .B(n12732), .C(n45), .Y(n4444) );
  NAND2X1 U53 ( .A(ram[7]), .B(n13035), .Y(n45) );
  OAI21X1 U54 ( .A(n13035), .B(n12726), .C(n46), .Y(n4445) );
  NAND2X1 U55 ( .A(ram[8]), .B(n13035), .Y(n46) );
  OAI21X1 U56 ( .A(n13035), .B(n12720), .C(n47), .Y(n4446) );
  NAND2X1 U57 ( .A(ram[9]), .B(n13035), .Y(n47) );
  OAI21X1 U58 ( .A(n13035), .B(n12714), .C(n48), .Y(n4447) );
  NAND2X1 U59 ( .A(ram[10]), .B(n13035), .Y(n48) );
  OAI21X1 U60 ( .A(n13035), .B(n12708), .C(n49), .Y(n4448) );
  NAND2X1 U61 ( .A(ram[11]), .B(n13035), .Y(n49) );
  OAI21X1 U62 ( .A(n13035), .B(n12702), .C(n50), .Y(n4449) );
  NAND2X1 U63 ( .A(ram[12]), .B(n13035), .Y(n50) );
  OAI21X1 U64 ( .A(n13035), .B(n12696), .C(n51), .Y(n4450) );
  NAND2X1 U65 ( .A(ram[13]), .B(n13035), .Y(n51) );
  OAI21X1 U66 ( .A(n13035), .B(n12692), .C(n52), .Y(n4451) );
  NAND2X1 U67 ( .A(ram[14]), .B(n13035), .Y(n52) );
  OAI21X1 U68 ( .A(n13035), .B(n12686), .C(n53), .Y(n4452) );
  NAND2X1 U69 ( .A(ram[15]), .B(n13035), .Y(n53) );
  OAI21X1 U71 ( .A(n13071), .B(n13034), .C(n56), .Y(n4453) );
  NAND2X1 U72 ( .A(ram[16]), .B(n13034), .Y(n56) );
  OAI21X1 U73 ( .A(n13070), .B(n13034), .C(n57), .Y(n4454) );
  NAND2X1 U74 ( .A(ram[17]), .B(n13034), .Y(n57) );
  OAI21X1 U75 ( .A(n12763), .B(n13034), .C(n58), .Y(n4455) );
  NAND2X1 U76 ( .A(ram[18]), .B(n13034), .Y(n58) );
  OAI21X1 U77 ( .A(n12757), .B(n13034), .C(n59), .Y(n4456) );
  NAND2X1 U78 ( .A(ram[19]), .B(n13034), .Y(n59) );
  OAI21X1 U79 ( .A(n12751), .B(n13034), .C(n60), .Y(n4457) );
  NAND2X1 U80 ( .A(ram[20]), .B(n13034), .Y(n60) );
  OAI21X1 U81 ( .A(n12745), .B(n13034), .C(n61), .Y(n4458) );
  NAND2X1 U82 ( .A(ram[21]), .B(n13034), .Y(n61) );
  OAI21X1 U83 ( .A(n12739), .B(n13034), .C(n62), .Y(n4459) );
  NAND2X1 U84 ( .A(ram[22]), .B(n13034), .Y(n62) );
  OAI21X1 U85 ( .A(n12733), .B(n13034), .C(n63), .Y(n4460) );
  NAND2X1 U86 ( .A(ram[23]), .B(n13034), .Y(n63) );
  OAI21X1 U87 ( .A(n12727), .B(n13034), .C(n64), .Y(n4461) );
  NAND2X1 U88 ( .A(ram[24]), .B(n13034), .Y(n64) );
  OAI21X1 U89 ( .A(n12721), .B(n13034), .C(n65), .Y(n4462) );
  NAND2X1 U90 ( .A(ram[25]), .B(n13034), .Y(n65) );
  OAI21X1 U91 ( .A(n12715), .B(n13034), .C(n66), .Y(n4463) );
  NAND2X1 U92 ( .A(ram[26]), .B(n13034), .Y(n66) );
  OAI21X1 U93 ( .A(n12709), .B(n13034), .C(n67), .Y(n4464) );
  NAND2X1 U94 ( .A(ram[27]), .B(n13034), .Y(n67) );
  OAI21X1 U95 ( .A(n12703), .B(n13034), .C(n68), .Y(n4465) );
  NAND2X1 U96 ( .A(ram[28]), .B(n13034), .Y(n68) );
  OAI21X1 U97 ( .A(n12697), .B(n13034), .C(n69), .Y(n4466) );
  NAND2X1 U98 ( .A(ram[29]), .B(n13034), .Y(n69) );
  OAI21X1 U99 ( .A(n13057), .B(n13034), .C(n70), .Y(n4467) );
  NAND2X1 U100 ( .A(ram[30]), .B(n13034), .Y(n70) );
  OAI21X1 U101 ( .A(n13056), .B(n13034), .C(n71), .Y(n4468) );
  NAND2X1 U102 ( .A(ram[31]), .B(n13034), .Y(n71) );
  OAI21X1 U104 ( .A(n13071), .B(n13033), .C(n74), .Y(n4469) );
  NAND2X1 U105 ( .A(ram[32]), .B(n13033), .Y(n74) );
  OAI21X1 U106 ( .A(n13070), .B(n13033), .C(n75), .Y(n4470) );
  NAND2X1 U107 ( .A(ram[33]), .B(n13033), .Y(n75) );
  OAI21X1 U108 ( .A(n12762), .B(n13033), .C(n76), .Y(n4471) );
  NAND2X1 U109 ( .A(ram[34]), .B(n13033), .Y(n76) );
  OAI21X1 U110 ( .A(n12756), .B(n13033), .C(n77), .Y(n4472) );
  NAND2X1 U111 ( .A(ram[35]), .B(n13033), .Y(n77) );
  OAI21X1 U112 ( .A(n12750), .B(n13033), .C(n78), .Y(n4473) );
  NAND2X1 U113 ( .A(ram[36]), .B(n13033), .Y(n78) );
  OAI21X1 U114 ( .A(n12744), .B(n13033), .C(n79), .Y(n4474) );
  NAND2X1 U115 ( .A(ram[37]), .B(n13033), .Y(n79) );
  OAI21X1 U116 ( .A(n12738), .B(n13033), .C(n80), .Y(n4475) );
  NAND2X1 U117 ( .A(ram[38]), .B(n13033), .Y(n80) );
  OAI21X1 U118 ( .A(n12732), .B(n13033), .C(n81), .Y(n4476) );
  NAND2X1 U119 ( .A(ram[39]), .B(n13033), .Y(n81) );
  OAI21X1 U120 ( .A(n12726), .B(n13033), .C(n82), .Y(n4477) );
  NAND2X1 U121 ( .A(ram[40]), .B(n13033), .Y(n82) );
  OAI21X1 U122 ( .A(n12720), .B(n13033), .C(n83), .Y(n4478) );
  NAND2X1 U123 ( .A(ram[41]), .B(n13033), .Y(n83) );
  OAI21X1 U124 ( .A(n12714), .B(n13033), .C(n84), .Y(n4479) );
  NAND2X1 U125 ( .A(ram[42]), .B(n13033), .Y(n84) );
  OAI21X1 U126 ( .A(n12708), .B(n13033), .C(n85), .Y(n4480) );
  NAND2X1 U127 ( .A(ram[43]), .B(n13033), .Y(n85) );
  OAI21X1 U128 ( .A(n12702), .B(n13033), .C(n86), .Y(n4481) );
  NAND2X1 U129 ( .A(ram[44]), .B(n13033), .Y(n86) );
  OAI21X1 U130 ( .A(n12696), .B(n13033), .C(n87), .Y(n4482) );
  NAND2X1 U131 ( .A(ram[45]), .B(n13033), .Y(n87) );
  OAI21X1 U132 ( .A(n13057), .B(n13033), .C(n88), .Y(n4483) );
  NAND2X1 U133 ( .A(ram[46]), .B(n13033), .Y(n88) );
  OAI21X1 U134 ( .A(n13056), .B(n13033), .C(n89), .Y(n4484) );
  NAND2X1 U135 ( .A(ram[47]), .B(n13033), .Y(n89) );
  OAI21X1 U137 ( .A(n13071), .B(n13032), .C(n92), .Y(n4485) );
  NAND2X1 U138 ( .A(ram[48]), .B(n13032), .Y(n92) );
  OAI21X1 U139 ( .A(n13070), .B(n13032), .C(n93), .Y(n4486) );
  NAND2X1 U140 ( .A(ram[49]), .B(n13032), .Y(n93) );
  OAI21X1 U141 ( .A(n12763), .B(n13032), .C(n94), .Y(n4487) );
  NAND2X1 U142 ( .A(ram[50]), .B(n13032), .Y(n94) );
  OAI21X1 U143 ( .A(n12757), .B(n13032), .C(n95), .Y(n4488) );
  NAND2X1 U144 ( .A(ram[51]), .B(n13032), .Y(n95) );
  OAI21X1 U145 ( .A(n12751), .B(n13032), .C(n96), .Y(n4489) );
  NAND2X1 U146 ( .A(ram[52]), .B(n13032), .Y(n96) );
  OAI21X1 U147 ( .A(n12745), .B(n13032), .C(n97), .Y(n4490) );
  NAND2X1 U148 ( .A(ram[53]), .B(n13032), .Y(n97) );
  OAI21X1 U149 ( .A(n12739), .B(n13032), .C(n98), .Y(n4491) );
  NAND2X1 U150 ( .A(ram[54]), .B(n13032), .Y(n98) );
  OAI21X1 U151 ( .A(n12733), .B(n13032), .C(n99), .Y(n4492) );
  NAND2X1 U152 ( .A(ram[55]), .B(n13032), .Y(n99) );
  OAI21X1 U153 ( .A(n12727), .B(n13032), .C(n100), .Y(n4493) );
  NAND2X1 U154 ( .A(ram[56]), .B(n13032), .Y(n100) );
  OAI21X1 U155 ( .A(n12721), .B(n13032), .C(n101), .Y(n4494) );
  NAND2X1 U156 ( .A(ram[57]), .B(n13032), .Y(n101) );
  OAI21X1 U157 ( .A(n12715), .B(n13032), .C(n102), .Y(n4495) );
  NAND2X1 U158 ( .A(ram[58]), .B(n13032), .Y(n102) );
  OAI21X1 U159 ( .A(n12709), .B(n13032), .C(n103), .Y(n4496) );
  NAND2X1 U160 ( .A(ram[59]), .B(n13032), .Y(n103) );
  OAI21X1 U161 ( .A(n12703), .B(n13032), .C(n104), .Y(n4497) );
  NAND2X1 U162 ( .A(ram[60]), .B(n13032), .Y(n104) );
  OAI21X1 U163 ( .A(n12697), .B(n13032), .C(n105), .Y(n4498) );
  NAND2X1 U164 ( .A(ram[61]), .B(n13032), .Y(n105) );
  OAI21X1 U165 ( .A(n13057), .B(n13032), .C(n106), .Y(n4499) );
  NAND2X1 U166 ( .A(ram[62]), .B(n13032), .Y(n106) );
  OAI21X1 U167 ( .A(n13056), .B(n13032), .C(n107), .Y(n4500) );
  NAND2X1 U168 ( .A(ram[63]), .B(n13032), .Y(n107) );
  OAI21X1 U170 ( .A(n13071), .B(n13031), .C(n110), .Y(n4501) );
  NAND2X1 U171 ( .A(ram[64]), .B(n13031), .Y(n110) );
  OAI21X1 U172 ( .A(n13070), .B(n13031), .C(n111), .Y(n4502) );
  NAND2X1 U173 ( .A(ram[65]), .B(n13031), .Y(n111) );
  OAI21X1 U174 ( .A(n13069), .B(n13031), .C(n112), .Y(n4503) );
  NAND2X1 U175 ( .A(ram[66]), .B(n13031), .Y(n112) );
  OAI21X1 U176 ( .A(n13068), .B(n13031), .C(n113), .Y(n4504) );
  NAND2X1 U177 ( .A(ram[67]), .B(n13031), .Y(n113) );
  OAI21X1 U178 ( .A(n13067), .B(n13031), .C(n114), .Y(n4505) );
  NAND2X1 U179 ( .A(ram[68]), .B(n13031), .Y(n114) );
  OAI21X1 U180 ( .A(n13066), .B(n13031), .C(n115), .Y(n4506) );
  NAND2X1 U181 ( .A(ram[69]), .B(n13031), .Y(n115) );
  OAI21X1 U182 ( .A(n13065), .B(n13031), .C(n116), .Y(n4507) );
  NAND2X1 U183 ( .A(ram[70]), .B(n13031), .Y(n116) );
  OAI21X1 U184 ( .A(n13064), .B(n13031), .C(n117), .Y(n4508) );
  NAND2X1 U185 ( .A(ram[71]), .B(n13031), .Y(n117) );
  OAI21X1 U186 ( .A(n13063), .B(n13031), .C(n118), .Y(n4509) );
  NAND2X1 U187 ( .A(ram[72]), .B(n13031), .Y(n118) );
  OAI21X1 U188 ( .A(n13062), .B(n13031), .C(n119), .Y(n4510) );
  NAND2X1 U189 ( .A(ram[73]), .B(n13031), .Y(n119) );
  OAI21X1 U190 ( .A(n13061), .B(n13031), .C(n120), .Y(n4511) );
  NAND2X1 U191 ( .A(ram[74]), .B(n13031), .Y(n120) );
  OAI21X1 U192 ( .A(n13060), .B(n13031), .C(n121), .Y(n4512) );
  NAND2X1 U193 ( .A(ram[75]), .B(n13031), .Y(n121) );
  OAI21X1 U194 ( .A(n13059), .B(n13031), .C(n122), .Y(n4513) );
  NAND2X1 U195 ( .A(ram[76]), .B(n13031), .Y(n122) );
  OAI21X1 U196 ( .A(n13058), .B(n13031), .C(n123), .Y(n4514) );
  NAND2X1 U197 ( .A(ram[77]), .B(n13031), .Y(n123) );
  OAI21X1 U198 ( .A(n13057), .B(n13031), .C(n124), .Y(n4515) );
  NAND2X1 U199 ( .A(ram[78]), .B(n13031), .Y(n124) );
  OAI21X1 U200 ( .A(n13056), .B(n13031), .C(n125), .Y(n4516) );
  NAND2X1 U201 ( .A(ram[79]), .B(n13031), .Y(n125) );
  OAI21X1 U203 ( .A(n13071), .B(n13030), .C(n128), .Y(n4517) );
  NAND2X1 U204 ( .A(ram[80]), .B(n13030), .Y(n128) );
  OAI21X1 U205 ( .A(n13070), .B(n13030), .C(n129), .Y(n4518) );
  NAND2X1 U206 ( .A(ram[81]), .B(n13030), .Y(n129) );
  OAI21X1 U207 ( .A(n13069), .B(n13030), .C(n130), .Y(n4519) );
  NAND2X1 U208 ( .A(ram[82]), .B(n13030), .Y(n130) );
  OAI21X1 U209 ( .A(n13068), .B(n13030), .C(n131), .Y(n4520) );
  NAND2X1 U210 ( .A(ram[83]), .B(n13030), .Y(n131) );
  OAI21X1 U211 ( .A(n13067), .B(n13030), .C(n132), .Y(n4521) );
  NAND2X1 U212 ( .A(ram[84]), .B(n13030), .Y(n132) );
  OAI21X1 U213 ( .A(n13066), .B(n13030), .C(n133), .Y(n4522) );
  NAND2X1 U214 ( .A(ram[85]), .B(n13030), .Y(n133) );
  OAI21X1 U215 ( .A(n13065), .B(n13030), .C(n134), .Y(n4523) );
  NAND2X1 U216 ( .A(ram[86]), .B(n13030), .Y(n134) );
  OAI21X1 U217 ( .A(n13064), .B(n13030), .C(n135), .Y(n4524) );
  NAND2X1 U218 ( .A(ram[87]), .B(n13030), .Y(n135) );
  OAI21X1 U219 ( .A(n13063), .B(n13030), .C(n136), .Y(n4525) );
  NAND2X1 U220 ( .A(ram[88]), .B(n13030), .Y(n136) );
  OAI21X1 U221 ( .A(n13062), .B(n13030), .C(n137), .Y(n4526) );
  NAND2X1 U222 ( .A(ram[89]), .B(n13030), .Y(n137) );
  OAI21X1 U223 ( .A(n13061), .B(n13030), .C(n138), .Y(n4527) );
  NAND2X1 U224 ( .A(ram[90]), .B(n13030), .Y(n138) );
  OAI21X1 U225 ( .A(n13060), .B(n13030), .C(n139), .Y(n4528) );
  NAND2X1 U226 ( .A(ram[91]), .B(n13030), .Y(n139) );
  OAI21X1 U227 ( .A(n13059), .B(n13030), .C(n140), .Y(n4529) );
  NAND2X1 U228 ( .A(ram[92]), .B(n13030), .Y(n140) );
  OAI21X1 U229 ( .A(n13058), .B(n13030), .C(n141), .Y(n4530) );
  NAND2X1 U230 ( .A(ram[93]), .B(n13030), .Y(n141) );
  OAI21X1 U231 ( .A(n13057), .B(n13030), .C(n142), .Y(n4531) );
  NAND2X1 U232 ( .A(ram[94]), .B(n13030), .Y(n142) );
  OAI21X1 U233 ( .A(n13056), .B(n13030), .C(n143), .Y(n4532) );
  NAND2X1 U234 ( .A(ram[95]), .B(n13030), .Y(n143) );
  OAI21X1 U236 ( .A(n13071), .B(n13029), .C(n146), .Y(n4533) );
  NAND2X1 U237 ( .A(ram[96]), .B(n13029), .Y(n146) );
  OAI21X1 U238 ( .A(n13070), .B(n13029), .C(n147), .Y(n4534) );
  NAND2X1 U239 ( .A(ram[97]), .B(n13029), .Y(n147) );
  OAI21X1 U240 ( .A(n13069), .B(n13029), .C(n148), .Y(n4535) );
  NAND2X1 U241 ( .A(ram[98]), .B(n13029), .Y(n148) );
  OAI21X1 U242 ( .A(n13068), .B(n13029), .C(n149), .Y(n4536) );
  NAND2X1 U243 ( .A(ram[99]), .B(n13029), .Y(n149) );
  OAI21X1 U244 ( .A(n13067), .B(n13029), .C(n150), .Y(n4537) );
  NAND2X1 U245 ( .A(ram[100]), .B(n13029), .Y(n150) );
  OAI21X1 U246 ( .A(n13066), .B(n13029), .C(n151), .Y(n4538) );
  NAND2X1 U247 ( .A(ram[101]), .B(n13029), .Y(n151) );
  OAI21X1 U248 ( .A(n13065), .B(n13029), .C(n152), .Y(n4539) );
  NAND2X1 U249 ( .A(ram[102]), .B(n13029), .Y(n152) );
  OAI21X1 U250 ( .A(n13064), .B(n13029), .C(n153), .Y(n4540) );
  NAND2X1 U251 ( .A(ram[103]), .B(n13029), .Y(n153) );
  OAI21X1 U252 ( .A(n13063), .B(n13029), .C(n154), .Y(n4541) );
  NAND2X1 U253 ( .A(ram[104]), .B(n13029), .Y(n154) );
  OAI21X1 U254 ( .A(n13062), .B(n13029), .C(n155), .Y(n4542) );
  NAND2X1 U255 ( .A(ram[105]), .B(n13029), .Y(n155) );
  OAI21X1 U256 ( .A(n13061), .B(n13029), .C(n156), .Y(n4543) );
  NAND2X1 U257 ( .A(ram[106]), .B(n13029), .Y(n156) );
  OAI21X1 U258 ( .A(n13060), .B(n13029), .C(n157), .Y(n4544) );
  NAND2X1 U259 ( .A(ram[107]), .B(n13029), .Y(n157) );
  OAI21X1 U260 ( .A(n13059), .B(n13029), .C(n158), .Y(n4545) );
  NAND2X1 U261 ( .A(ram[108]), .B(n13029), .Y(n158) );
  OAI21X1 U262 ( .A(n13058), .B(n13029), .C(n159), .Y(n4546) );
  NAND2X1 U263 ( .A(ram[109]), .B(n13029), .Y(n159) );
  OAI21X1 U264 ( .A(n13057), .B(n13029), .C(n160), .Y(n4547) );
  NAND2X1 U265 ( .A(ram[110]), .B(n13029), .Y(n160) );
  OAI21X1 U266 ( .A(n13056), .B(n13029), .C(n161), .Y(n4548) );
  NAND2X1 U267 ( .A(ram[111]), .B(n13029), .Y(n161) );
  OAI21X1 U269 ( .A(n13071), .B(n13028), .C(n164), .Y(n4549) );
  NAND2X1 U270 ( .A(ram[112]), .B(n13028), .Y(n164) );
  OAI21X1 U271 ( .A(n13070), .B(n13028), .C(n165), .Y(n4550) );
  NAND2X1 U272 ( .A(ram[113]), .B(n13028), .Y(n165) );
  OAI21X1 U273 ( .A(n13069), .B(n13028), .C(n166), .Y(n4551) );
  NAND2X1 U274 ( .A(ram[114]), .B(n13028), .Y(n166) );
  OAI21X1 U275 ( .A(n13068), .B(n13028), .C(n167), .Y(n4552) );
  NAND2X1 U276 ( .A(ram[115]), .B(n13028), .Y(n167) );
  OAI21X1 U277 ( .A(n13067), .B(n13028), .C(n168), .Y(n4553) );
  NAND2X1 U278 ( .A(ram[116]), .B(n13028), .Y(n168) );
  OAI21X1 U279 ( .A(n13066), .B(n13028), .C(n169), .Y(n4554) );
  NAND2X1 U280 ( .A(ram[117]), .B(n13028), .Y(n169) );
  OAI21X1 U281 ( .A(n13065), .B(n13028), .C(n170), .Y(n4555) );
  NAND2X1 U282 ( .A(ram[118]), .B(n13028), .Y(n170) );
  OAI21X1 U283 ( .A(n13064), .B(n13028), .C(n171), .Y(n4556) );
  NAND2X1 U284 ( .A(ram[119]), .B(n13028), .Y(n171) );
  OAI21X1 U285 ( .A(n13063), .B(n13028), .C(n172), .Y(n4557) );
  NAND2X1 U286 ( .A(ram[120]), .B(n13028), .Y(n172) );
  OAI21X1 U287 ( .A(n13062), .B(n13028), .C(n173), .Y(n4558) );
  NAND2X1 U288 ( .A(ram[121]), .B(n13028), .Y(n173) );
  OAI21X1 U289 ( .A(n13061), .B(n13028), .C(n174), .Y(n4559) );
  NAND2X1 U290 ( .A(ram[122]), .B(n13028), .Y(n174) );
  OAI21X1 U291 ( .A(n13060), .B(n13028), .C(n175), .Y(n4560) );
  NAND2X1 U292 ( .A(ram[123]), .B(n13028), .Y(n175) );
  OAI21X1 U293 ( .A(n13059), .B(n13028), .C(n176), .Y(n4561) );
  NAND2X1 U294 ( .A(ram[124]), .B(n13028), .Y(n176) );
  OAI21X1 U295 ( .A(n13058), .B(n13028), .C(n177), .Y(n4562) );
  NAND2X1 U296 ( .A(ram[125]), .B(n13028), .Y(n177) );
  OAI21X1 U297 ( .A(n13057), .B(n13028), .C(n178), .Y(n4563) );
  NAND2X1 U298 ( .A(ram[126]), .B(n13028), .Y(n178) );
  OAI21X1 U299 ( .A(n13056), .B(n13028), .C(n179), .Y(n4564) );
  NAND2X1 U300 ( .A(ram[127]), .B(n13028), .Y(n179) );
  OAI21X1 U302 ( .A(n13071), .B(n13027), .C(n182), .Y(n4565) );
  NAND2X1 U303 ( .A(ram[128]), .B(n13027), .Y(n182) );
  OAI21X1 U304 ( .A(n13070), .B(n13027), .C(n183), .Y(n4566) );
  NAND2X1 U305 ( .A(ram[129]), .B(n13027), .Y(n183) );
  OAI21X1 U306 ( .A(n13069), .B(n13027), .C(n184), .Y(n4567) );
  NAND2X1 U307 ( .A(ram[130]), .B(n13027), .Y(n184) );
  OAI21X1 U308 ( .A(n13068), .B(n13027), .C(n185), .Y(n4568) );
  NAND2X1 U309 ( .A(ram[131]), .B(n13027), .Y(n185) );
  OAI21X1 U310 ( .A(n13067), .B(n13027), .C(n186), .Y(n4569) );
  NAND2X1 U311 ( .A(ram[132]), .B(n13027), .Y(n186) );
  OAI21X1 U312 ( .A(n13066), .B(n13027), .C(n187), .Y(n4570) );
  NAND2X1 U313 ( .A(ram[133]), .B(n13027), .Y(n187) );
  OAI21X1 U314 ( .A(n13065), .B(n13027), .C(n188), .Y(n4571) );
  NAND2X1 U315 ( .A(ram[134]), .B(n13027), .Y(n188) );
  OAI21X1 U316 ( .A(n13064), .B(n13027), .C(n189), .Y(n4572) );
  NAND2X1 U317 ( .A(ram[135]), .B(n13027), .Y(n189) );
  OAI21X1 U318 ( .A(n13063), .B(n13027), .C(n190), .Y(n4573) );
  NAND2X1 U319 ( .A(ram[136]), .B(n13027), .Y(n190) );
  OAI21X1 U320 ( .A(n13062), .B(n13027), .C(n191), .Y(n4574) );
  NAND2X1 U321 ( .A(ram[137]), .B(n13027), .Y(n191) );
  OAI21X1 U322 ( .A(n13061), .B(n13027), .C(n192), .Y(n4575) );
  NAND2X1 U323 ( .A(ram[138]), .B(n13027), .Y(n192) );
  OAI21X1 U324 ( .A(n13060), .B(n13027), .C(n193), .Y(n4576) );
  NAND2X1 U325 ( .A(ram[139]), .B(n13027), .Y(n193) );
  OAI21X1 U326 ( .A(n13059), .B(n13027), .C(n194), .Y(n4577) );
  NAND2X1 U327 ( .A(ram[140]), .B(n13027), .Y(n194) );
  OAI21X1 U328 ( .A(n13058), .B(n13027), .C(n195), .Y(n4578) );
  NAND2X1 U329 ( .A(ram[141]), .B(n13027), .Y(n195) );
  OAI21X1 U330 ( .A(n13057), .B(n13027), .C(n196), .Y(n4579) );
  NAND2X1 U331 ( .A(ram[142]), .B(n13027), .Y(n196) );
  OAI21X1 U332 ( .A(n13056), .B(n13027), .C(n197), .Y(n4580) );
  NAND2X1 U333 ( .A(ram[143]), .B(n13027), .Y(n197) );
  OAI21X1 U335 ( .A(n13071), .B(n13026), .C(n200), .Y(n4581) );
  NAND2X1 U336 ( .A(ram[144]), .B(n13026), .Y(n200) );
  OAI21X1 U337 ( .A(n13070), .B(n13026), .C(n201), .Y(n4582) );
  NAND2X1 U338 ( .A(ram[145]), .B(n13026), .Y(n201) );
  OAI21X1 U339 ( .A(n13069), .B(n13026), .C(n202), .Y(n4583) );
  NAND2X1 U340 ( .A(ram[146]), .B(n13026), .Y(n202) );
  OAI21X1 U341 ( .A(n13068), .B(n13026), .C(n203), .Y(n4584) );
  NAND2X1 U342 ( .A(ram[147]), .B(n13026), .Y(n203) );
  OAI21X1 U343 ( .A(n13067), .B(n13026), .C(n204), .Y(n4585) );
  NAND2X1 U344 ( .A(ram[148]), .B(n13026), .Y(n204) );
  OAI21X1 U345 ( .A(n13066), .B(n13026), .C(n205), .Y(n4586) );
  NAND2X1 U346 ( .A(ram[149]), .B(n13026), .Y(n205) );
  OAI21X1 U347 ( .A(n13065), .B(n13026), .C(n206), .Y(n4587) );
  NAND2X1 U348 ( .A(ram[150]), .B(n13026), .Y(n206) );
  OAI21X1 U349 ( .A(n13064), .B(n13026), .C(n207), .Y(n4588) );
  NAND2X1 U350 ( .A(ram[151]), .B(n13026), .Y(n207) );
  OAI21X1 U351 ( .A(n13063), .B(n13026), .C(n208), .Y(n4589) );
  NAND2X1 U352 ( .A(ram[152]), .B(n13026), .Y(n208) );
  OAI21X1 U353 ( .A(n13062), .B(n13026), .C(n209), .Y(n4590) );
  NAND2X1 U354 ( .A(ram[153]), .B(n13026), .Y(n209) );
  OAI21X1 U355 ( .A(n13061), .B(n13026), .C(n210), .Y(n4591) );
  NAND2X1 U356 ( .A(ram[154]), .B(n13026), .Y(n210) );
  OAI21X1 U357 ( .A(n13060), .B(n13026), .C(n211), .Y(n4592) );
  NAND2X1 U358 ( .A(ram[155]), .B(n13026), .Y(n211) );
  OAI21X1 U359 ( .A(n13059), .B(n13026), .C(n212), .Y(n4593) );
  NAND2X1 U360 ( .A(ram[156]), .B(n13026), .Y(n212) );
  OAI21X1 U361 ( .A(n13058), .B(n13026), .C(n213), .Y(n4594) );
  NAND2X1 U362 ( .A(ram[157]), .B(n13026), .Y(n213) );
  OAI21X1 U363 ( .A(n13057), .B(n13026), .C(n214), .Y(n4595) );
  NAND2X1 U364 ( .A(ram[158]), .B(n13026), .Y(n214) );
  OAI21X1 U365 ( .A(n13056), .B(n13026), .C(n215), .Y(n4596) );
  NAND2X1 U366 ( .A(ram[159]), .B(n13026), .Y(n215) );
  OAI21X1 U368 ( .A(n12777), .B(n13025), .C(n218), .Y(n4597) );
  NAND2X1 U369 ( .A(ram[160]), .B(n13025), .Y(n218) );
  OAI21X1 U370 ( .A(n12771), .B(n13025), .C(n219), .Y(n4598) );
  NAND2X1 U371 ( .A(ram[161]), .B(n13025), .Y(n219) );
  OAI21X1 U372 ( .A(n12764), .B(n13025), .C(n220), .Y(n4599) );
  NAND2X1 U373 ( .A(ram[162]), .B(n13025), .Y(n220) );
  OAI21X1 U374 ( .A(n12758), .B(n13025), .C(n221), .Y(n4600) );
  NAND2X1 U375 ( .A(ram[163]), .B(n13025), .Y(n221) );
  OAI21X1 U376 ( .A(n12752), .B(n13025), .C(n222), .Y(n4601) );
  NAND2X1 U377 ( .A(ram[164]), .B(n13025), .Y(n222) );
  OAI21X1 U378 ( .A(n12746), .B(n13025), .C(n223), .Y(n4602) );
  NAND2X1 U379 ( .A(ram[165]), .B(n13025), .Y(n223) );
  OAI21X1 U380 ( .A(n12740), .B(n13025), .C(n224), .Y(n4603) );
  NAND2X1 U381 ( .A(ram[166]), .B(n13025), .Y(n224) );
  OAI21X1 U382 ( .A(n12734), .B(n13025), .C(n225), .Y(n4604) );
  NAND2X1 U383 ( .A(ram[167]), .B(n13025), .Y(n225) );
  OAI21X1 U384 ( .A(n12728), .B(n13025), .C(n226), .Y(n4605) );
  NAND2X1 U385 ( .A(ram[168]), .B(n13025), .Y(n226) );
  OAI21X1 U386 ( .A(n12722), .B(n13025), .C(n227), .Y(n4606) );
  NAND2X1 U387 ( .A(ram[169]), .B(n13025), .Y(n227) );
  OAI21X1 U388 ( .A(n12716), .B(n13025), .C(n228), .Y(n4607) );
  NAND2X1 U389 ( .A(ram[170]), .B(n13025), .Y(n228) );
  OAI21X1 U390 ( .A(n12710), .B(n13025), .C(n229), .Y(n4608) );
  NAND2X1 U391 ( .A(ram[171]), .B(n13025), .Y(n229) );
  OAI21X1 U392 ( .A(n12704), .B(n13025), .C(n230), .Y(n4609) );
  NAND2X1 U393 ( .A(ram[172]), .B(n13025), .Y(n230) );
  OAI21X1 U394 ( .A(n12698), .B(n13025), .C(n231), .Y(n4610) );
  NAND2X1 U395 ( .A(ram[173]), .B(n13025), .Y(n231) );
  OAI21X1 U396 ( .A(n12693), .B(n13025), .C(n232), .Y(n4611) );
  NAND2X1 U397 ( .A(ram[174]), .B(n13025), .Y(n232) );
  OAI21X1 U398 ( .A(n12687), .B(n13025), .C(n233), .Y(n4612) );
  NAND2X1 U399 ( .A(ram[175]), .B(n13025), .Y(n233) );
  OAI21X1 U401 ( .A(n12775), .B(n13024), .C(n236), .Y(n4613) );
  NAND2X1 U402 ( .A(ram[176]), .B(n13024), .Y(n236) );
  OAI21X1 U403 ( .A(n12769), .B(n13024), .C(n237), .Y(n4614) );
  NAND2X1 U404 ( .A(ram[177]), .B(n13024), .Y(n237) );
  OAI21X1 U405 ( .A(n12762), .B(n13024), .C(n238), .Y(n4615) );
  NAND2X1 U406 ( .A(ram[178]), .B(n13024), .Y(n238) );
  OAI21X1 U407 ( .A(n12756), .B(n13024), .C(n239), .Y(n4616) );
  NAND2X1 U408 ( .A(ram[179]), .B(n13024), .Y(n239) );
  OAI21X1 U409 ( .A(n12750), .B(n13024), .C(n240), .Y(n4617) );
  NAND2X1 U410 ( .A(ram[180]), .B(n13024), .Y(n240) );
  OAI21X1 U411 ( .A(n12744), .B(n13024), .C(n241), .Y(n4618) );
  NAND2X1 U412 ( .A(ram[181]), .B(n13024), .Y(n241) );
  OAI21X1 U413 ( .A(n12738), .B(n13024), .C(n242), .Y(n4619) );
  NAND2X1 U414 ( .A(ram[182]), .B(n13024), .Y(n242) );
  OAI21X1 U415 ( .A(n12732), .B(n13024), .C(n243), .Y(n4620) );
  NAND2X1 U416 ( .A(ram[183]), .B(n13024), .Y(n243) );
  OAI21X1 U417 ( .A(n12726), .B(n13024), .C(n244), .Y(n4621) );
  NAND2X1 U418 ( .A(ram[184]), .B(n13024), .Y(n244) );
  OAI21X1 U419 ( .A(n12720), .B(n13024), .C(n245), .Y(n4622) );
  NAND2X1 U420 ( .A(ram[185]), .B(n13024), .Y(n245) );
  OAI21X1 U421 ( .A(n12714), .B(n13024), .C(n246), .Y(n4623) );
  NAND2X1 U422 ( .A(ram[186]), .B(n13024), .Y(n246) );
  OAI21X1 U423 ( .A(n12708), .B(n13024), .C(n247), .Y(n4624) );
  NAND2X1 U424 ( .A(ram[187]), .B(n13024), .Y(n247) );
  OAI21X1 U425 ( .A(n12702), .B(n13024), .C(n248), .Y(n4625) );
  NAND2X1 U426 ( .A(ram[188]), .B(n13024), .Y(n248) );
  OAI21X1 U427 ( .A(n12696), .B(n13024), .C(n249), .Y(n4626) );
  NAND2X1 U428 ( .A(ram[189]), .B(n13024), .Y(n249) );
  OAI21X1 U429 ( .A(n12691), .B(n13024), .C(n250), .Y(n4627) );
  NAND2X1 U430 ( .A(ram[190]), .B(n13024), .Y(n250) );
  OAI21X1 U431 ( .A(n12685), .B(n13024), .C(n251), .Y(n4628) );
  NAND2X1 U432 ( .A(ram[191]), .B(n13024), .Y(n251) );
  OAI21X1 U434 ( .A(n12774), .B(n13023), .C(n254), .Y(n4629) );
  NAND2X1 U435 ( .A(ram[192]), .B(n13023), .Y(n254) );
  OAI21X1 U436 ( .A(n12768), .B(n13023), .C(n255), .Y(n4630) );
  NAND2X1 U437 ( .A(ram[193]), .B(n13023), .Y(n255) );
  OAI21X1 U438 ( .A(n12763), .B(n13023), .C(n256), .Y(n4631) );
  NAND2X1 U439 ( .A(ram[194]), .B(n13023), .Y(n256) );
  OAI21X1 U440 ( .A(n12757), .B(n13023), .C(n257), .Y(n4632) );
  NAND2X1 U441 ( .A(ram[195]), .B(n13023), .Y(n257) );
  OAI21X1 U442 ( .A(n12751), .B(n13023), .C(n258), .Y(n4633) );
  NAND2X1 U443 ( .A(ram[196]), .B(n13023), .Y(n258) );
  OAI21X1 U444 ( .A(n12745), .B(n13023), .C(n259), .Y(n4634) );
  NAND2X1 U445 ( .A(ram[197]), .B(n13023), .Y(n259) );
  OAI21X1 U446 ( .A(n12739), .B(n13023), .C(n260), .Y(n4635) );
  NAND2X1 U447 ( .A(ram[198]), .B(n13023), .Y(n260) );
  OAI21X1 U448 ( .A(n12733), .B(n13023), .C(n261), .Y(n4636) );
  NAND2X1 U449 ( .A(ram[199]), .B(n13023), .Y(n261) );
  OAI21X1 U450 ( .A(n12727), .B(n13023), .C(n262), .Y(n4637) );
  NAND2X1 U451 ( .A(ram[200]), .B(n13023), .Y(n262) );
  OAI21X1 U452 ( .A(n12721), .B(n13023), .C(n263), .Y(n4638) );
  NAND2X1 U453 ( .A(ram[201]), .B(n13023), .Y(n263) );
  OAI21X1 U454 ( .A(n12715), .B(n13023), .C(n264), .Y(n4639) );
  NAND2X1 U455 ( .A(ram[202]), .B(n13023), .Y(n264) );
  OAI21X1 U456 ( .A(n12709), .B(n13023), .C(n265), .Y(n4640) );
  NAND2X1 U457 ( .A(ram[203]), .B(n13023), .Y(n265) );
  OAI21X1 U458 ( .A(n12703), .B(n13023), .C(n266), .Y(n4641) );
  NAND2X1 U459 ( .A(ram[204]), .B(n13023), .Y(n266) );
  OAI21X1 U460 ( .A(n12697), .B(n13023), .C(n267), .Y(n4642) );
  NAND2X1 U461 ( .A(ram[205]), .B(n13023), .Y(n267) );
  OAI21X1 U462 ( .A(n12690), .B(n13023), .C(n268), .Y(n4643) );
  NAND2X1 U463 ( .A(ram[206]), .B(n13023), .Y(n268) );
  OAI21X1 U464 ( .A(n12684), .B(n13023), .C(n269), .Y(n4644) );
  NAND2X1 U465 ( .A(ram[207]), .B(n13023), .Y(n269) );
  OAI21X1 U467 ( .A(n13071), .B(n13022), .C(n272), .Y(n4645) );
  NAND2X1 U468 ( .A(ram[208]), .B(n13022), .Y(n272) );
  OAI21X1 U469 ( .A(n13070), .B(n13022), .C(n273), .Y(n4646) );
  NAND2X1 U470 ( .A(ram[209]), .B(n13022), .Y(n273) );
  OAI21X1 U471 ( .A(n13069), .B(n13022), .C(n274), .Y(n4647) );
  NAND2X1 U472 ( .A(ram[210]), .B(n13022), .Y(n274) );
  OAI21X1 U473 ( .A(n13068), .B(n13022), .C(n275), .Y(n4648) );
  NAND2X1 U474 ( .A(ram[211]), .B(n13022), .Y(n275) );
  OAI21X1 U475 ( .A(n13067), .B(n13022), .C(n276), .Y(n4649) );
  NAND2X1 U476 ( .A(ram[212]), .B(n13022), .Y(n276) );
  OAI21X1 U477 ( .A(n13066), .B(n13022), .C(n277), .Y(n4650) );
  NAND2X1 U478 ( .A(ram[213]), .B(n13022), .Y(n277) );
  OAI21X1 U479 ( .A(n13065), .B(n13022), .C(n278), .Y(n4651) );
  NAND2X1 U480 ( .A(ram[214]), .B(n13022), .Y(n278) );
  OAI21X1 U481 ( .A(n13064), .B(n13022), .C(n279), .Y(n4652) );
  NAND2X1 U482 ( .A(ram[215]), .B(n13022), .Y(n279) );
  OAI21X1 U483 ( .A(n13063), .B(n13022), .C(n280), .Y(n4653) );
  NAND2X1 U484 ( .A(ram[216]), .B(n13022), .Y(n280) );
  OAI21X1 U485 ( .A(n13062), .B(n13022), .C(n281), .Y(n4654) );
  NAND2X1 U486 ( .A(ram[217]), .B(n13022), .Y(n281) );
  OAI21X1 U487 ( .A(n13061), .B(n13022), .C(n282), .Y(n4655) );
  NAND2X1 U488 ( .A(ram[218]), .B(n13022), .Y(n282) );
  OAI21X1 U489 ( .A(n13060), .B(n13022), .C(n283), .Y(n4656) );
  NAND2X1 U490 ( .A(ram[219]), .B(n13022), .Y(n283) );
  OAI21X1 U491 ( .A(n13059), .B(n13022), .C(n284), .Y(n4657) );
  NAND2X1 U492 ( .A(ram[220]), .B(n13022), .Y(n284) );
  OAI21X1 U493 ( .A(n13058), .B(n13022), .C(n285), .Y(n4658) );
  NAND2X1 U494 ( .A(ram[221]), .B(n13022), .Y(n285) );
  OAI21X1 U495 ( .A(n13057), .B(n13022), .C(n286), .Y(n4659) );
  NAND2X1 U496 ( .A(ram[222]), .B(n13022), .Y(n286) );
  OAI21X1 U497 ( .A(n13056), .B(n13022), .C(n287), .Y(n4660) );
  NAND2X1 U498 ( .A(ram[223]), .B(n13022), .Y(n287) );
  OAI21X1 U500 ( .A(n13071), .B(n13021), .C(n290), .Y(n4661) );
  NAND2X1 U501 ( .A(ram[224]), .B(n13021), .Y(n290) );
  OAI21X1 U502 ( .A(n13070), .B(n13021), .C(n291), .Y(n4662) );
  NAND2X1 U503 ( .A(ram[225]), .B(n13021), .Y(n291) );
  OAI21X1 U504 ( .A(n13069), .B(n13021), .C(n292), .Y(n4663) );
  NAND2X1 U505 ( .A(ram[226]), .B(n13021), .Y(n292) );
  OAI21X1 U506 ( .A(n13068), .B(n13021), .C(n293), .Y(n4664) );
  NAND2X1 U507 ( .A(ram[227]), .B(n13021), .Y(n293) );
  OAI21X1 U508 ( .A(n13067), .B(n13021), .C(n294), .Y(n4665) );
  NAND2X1 U509 ( .A(ram[228]), .B(n13021), .Y(n294) );
  OAI21X1 U510 ( .A(n13066), .B(n13021), .C(n295), .Y(n4666) );
  NAND2X1 U511 ( .A(ram[229]), .B(n13021), .Y(n295) );
  OAI21X1 U512 ( .A(n13065), .B(n13021), .C(n296), .Y(n4667) );
  NAND2X1 U513 ( .A(ram[230]), .B(n13021), .Y(n296) );
  OAI21X1 U514 ( .A(n13064), .B(n13021), .C(n297), .Y(n4668) );
  NAND2X1 U515 ( .A(ram[231]), .B(n13021), .Y(n297) );
  OAI21X1 U516 ( .A(n13063), .B(n13021), .C(n298), .Y(n4669) );
  NAND2X1 U517 ( .A(ram[232]), .B(n13021), .Y(n298) );
  OAI21X1 U518 ( .A(n13062), .B(n13021), .C(n299), .Y(n4670) );
  NAND2X1 U519 ( .A(ram[233]), .B(n13021), .Y(n299) );
  OAI21X1 U520 ( .A(n13061), .B(n13021), .C(n300), .Y(n4671) );
  NAND2X1 U521 ( .A(ram[234]), .B(n13021), .Y(n300) );
  OAI21X1 U522 ( .A(n13060), .B(n13021), .C(n301), .Y(n4672) );
  NAND2X1 U523 ( .A(ram[235]), .B(n13021), .Y(n301) );
  OAI21X1 U524 ( .A(n13059), .B(n13021), .C(n302), .Y(n4673) );
  NAND2X1 U525 ( .A(ram[236]), .B(n13021), .Y(n302) );
  OAI21X1 U526 ( .A(n13058), .B(n13021), .C(n303), .Y(n4674) );
  NAND2X1 U527 ( .A(ram[237]), .B(n13021), .Y(n303) );
  OAI21X1 U528 ( .A(n13057), .B(n13021), .C(n304), .Y(n4675) );
  NAND2X1 U529 ( .A(ram[238]), .B(n13021), .Y(n304) );
  OAI21X1 U530 ( .A(n13056), .B(n13021), .C(n305), .Y(n4676) );
  NAND2X1 U531 ( .A(ram[239]), .B(n13021), .Y(n305) );
  OAI21X1 U533 ( .A(n13071), .B(n13020), .C(n308), .Y(n4677) );
  NAND2X1 U534 ( .A(ram[240]), .B(n13020), .Y(n308) );
  OAI21X1 U535 ( .A(n13070), .B(n13020), .C(n309), .Y(n4678) );
  NAND2X1 U536 ( .A(ram[241]), .B(n13020), .Y(n309) );
  OAI21X1 U537 ( .A(n13069), .B(n13020), .C(n310), .Y(n4679) );
  NAND2X1 U538 ( .A(ram[242]), .B(n13020), .Y(n310) );
  OAI21X1 U539 ( .A(n13068), .B(n13020), .C(n311), .Y(n4680) );
  NAND2X1 U540 ( .A(ram[243]), .B(n13020), .Y(n311) );
  OAI21X1 U541 ( .A(n13067), .B(n13020), .C(n312), .Y(n4681) );
  NAND2X1 U542 ( .A(ram[244]), .B(n13020), .Y(n312) );
  OAI21X1 U543 ( .A(n13066), .B(n13020), .C(n313), .Y(n4682) );
  NAND2X1 U544 ( .A(ram[245]), .B(n13020), .Y(n313) );
  OAI21X1 U545 ( .A(n13065), .B(n13020), .C(n314), .Y(n4683) );
  NAND2X1 U546 ( .A(ram[246]), .B(n13020), .Y(n314) );
  OAI21X1 U547 ( .A(n13064), .B(n13020), .C(n315), .Y(n4684) );
  NAND2X1 U548 ( .A(ram[247]), .B(n13020), .Y(n315) );
  OAI21X1 U549 ( .A(n13063), .B(n13020), .C(n316), .Y(n4685) );
  NAND2X1 U550 ( .A(ram[248]), .B(n13020), .Y(n316) );
  OAI21X1 U551 ( .A(n13062), .B(n13020), .C(n317), .Y(n4686) );
  NAND2X1 U552 ( .A(ram[249]), .B(n13020), .Y(n317) );
  OAI21X1 U553 ( .A(n13061), .B(n13020), .C(n318), .Y(n4687) );
  NAND2X1 U554 ( .A(ram[250]), .B(n13020), .Y(n318) );
  OAI21X1 U555 ( .A(n13060), .B(n13020), .C(n319), .Y(n4688) );
  NAND2X1 U556 ( .A(ram[251]), .B(n13020), .Y(n319) );
  OAI21X1 U557 ( .A(n13059), .B(n13020), .C(n320), .Y(n4689) );
  NAND2X1 U558 ( .A(ram[252]), .B(n13020), .Y(n320) );
  OAI21X1 U559 ( .A(n13058), .B(n13020), .C(n321), .Y(n4690) );
  NAND2X1 U560 ( .A(ram[253]), .B(n13020), .Y(n321) );
  OAI21X1 U561 ( .A(n13057), .B(n13020), .C(n322), .Y(n4691) );
  NAND2X1 U562 ( .A(ram[254]), .B(n13020), .Y(n322) );
  OAI21X1 U563 ( .A(n13056), .B(n13020), .C(n323), .Y(n4692) );
  NAND2X1 U564 ( .A(ram[255]), .B(n13020), .Y(n323) );
  NAND3X1 U566 ( .A(n326), .B(n327), .C(mem_write_en), .Y(n325) );
  OAI21X1 U567 ( .A(n13071), .B(n13019), .C(n329), .Y(n4693) );
  NAND2X1 U568 ( .A(ram[256]), .B(n13019), .Y(n329) );
  OAI21X1 U569 ( .A(n13070), .B(n13019), .C(n330), .Y(n4694) );
  NAND2X1 U570 ( .A(ram[257]), .B(n13019), .Y(n330) );
  OAI21X1 U571 ( .A(n13069), .B(n13019), .C(n331), .Y(n4695) );
  NAND2X1 U572 ( .A(ram[258]), .B(n13019), .Y(n331) );
  OAI21X1 U573 ( .A(n13068), .B(n13019), .C(n332), .Y(n4696) );
  NAND2X1 U574 ( .A(ram[259]), .B(n13019), .Y(n332) );
  OAI21X1 U575 ( .A(n13067), .B(n13019), .C(n333), .Y(n4697) );
  NAND2X1 U576 ( .A(ram[260]), .B(n13019), .Y(n333) );
  OAI21X1 U577 ( .A(n13066), .B(n13019), .C(n334), .Y(n4698) );
  NAND2X1 U578 ( .A(ram[261]), .B(n13019), .Y(n334) );
  OAI21X1 U579 ( .A(n13065), .B(n13019), .C(n335), .Y(n4699) );
  NAND2X1 U580 ( .A(ram[262]), .B(n13019), .Y(n335) );
  OAI21X1 U581 ( .A(n13064), .B(n13019), .C(n336), .Y(n4700) );
  NAND2X1 U582 ( .A(ram[263]), .B(n13019), .Y(n336) );
  OAI21X1 U583 ( .A(n13063), .B(n13019), .C(n337), .Y(n4701) );
  NAND2X1 U584 ( .A(ram[264]), .B(n13019), .Y(n337) );
  OAI21X1 U585 ( .A(n13062), .B(n13019), .C(n338), .Y(n4702) );
  NAND2X1 U586 ( .A(ram[265]), .B(n13019), .Y(n338) );
  OAI21X1 U587 ( .A(n13061), .B(n13019), .C(n339), .Y(n4703) );
  NAND2X1 U588 ( .A(ram[266]), .B(n13019), .Y(n339) );
  OAI21X1 U589 ( .A(n13060), .B(n13019), .C(n340), .Y(n4704) );
  NAND2X1 U590 ( .A(ram[267]), .B(n13019), .Y(n340) );
  OAI21X1 U591 ( .A(n13059), .B(n13019), .C(n341), .Y(n4705) );
  NAND2X1 U592 ( .A(ram[268]), .B(n13019), .Y(n341) );
  OAI21X1 U593 ( .A(n13058), .B(n13019), .C(n342), .Y(n4706) );
  NAND2X1 U594 ( .A(ram[269]), .B(n13019), .Y(n342) );
  OAI21X1 U595 ( .A(n13057), .B(n13019), .C(n343), .Y(n4707) );
  NAND2X1 U596 ( .A(ram[270]), .B(n13019), .Y(n343) );
  OAI21X1 U597 ( .A(n13056), .B(n13019), .C(n344), .Y(n4708) );
  NAND2X1 U598 ( .A(ram[271]), .B(n13019), .Y(n344) );
  OAI21X1 U600 ( .A(n13071), .B(n13018), .C(n346), .Y(n4709) );
  NAND2X1 U601 ( .A(ram[272]), .B(n13018), .Y(n346) );
  OAI21X1 U602 ( .A(n13070), .B(n13018), .C(n347), .Y(n4710) );
  NAND2X1 U603 ( .A(ram[273]), .B(n13018), .Y(n347) );
  OAI21X1 U604 ( .A(n13069), .B(n13018), .C(n348), .Y(n4711) );
  NAND2X1 U605 ( .A(ram[274]), .B(n13018), .Y(n348) );
  OAI21X1 U606 ( .A(n13068), .B(n13018), .C(n349), .Y(n4712) );
  NAND2X1 U607 ( .A(ram[275]), .B(n13018), .Y(n349) );
  OAI21X1 U608 ( .A(n13067), .B(n13018), .C(n350), .Y(n4713) );
  NAND2X1 U609 ( .A(ram[276]), .B(n13018), .Y(n350) );
  OAI21X1 U610 ( .A(n13066), .B(n13018), .C(n351), .Y(n4714) );
  NAND2X1 U611 ( .A(ram[277]), .B(n13018), .Y(n351) );
  OAI21X1 U612 ( .A(n13065), .B(n13018), .C(n352), .Y(n4715) );
  NAND2X1 U613 ( .A(ram[278]), .B(n13018), .Y(n352) );
  OAI21X1 U614 ( .A(n13064), .B(n13018), .C(n353), .Y(n4716) );
  NAND2X1 U615 ( .A(ram[279]), .B(n13018), .Y(n353) );
  OAI21X1 U616 ( .A(n13063), .B(n13018), .C(n354), .Y(n4717) );
  NAND2X1 U617 ( .A(ram[280]), .B(n13018), .Y(n354) );
  OAI21X1 U618 ( .A(n13062), .B(n13018), .C(n355), .Y(n4718) );
  NAND2X1 U619 ( .A(ram[281]), .B(n13018), .Y(n355) );
  OAI21X1 U620 ( .A(n13061), .B(n13018), .C(n356), .Y(n4719) );
  NAND2X1 U621 ( .A(ram[282]), .B(n13018), .Y(n356) );
  OAI21X1 U622 ( .A(n13060), .B(n13018), .C(n357), .Y(n4720) );
  NAND2X1 U623 ( .A(ram[283]), .B(n13018), .Y(n357) );
  OAI21X1 U624 ( .A(n13059), .B(n13018), .C(n358), .Y(n4721) );
  NAND2X1 U625 ( .A(ram[284]), .B(n13018), .Y(n358) );
  OAI21X1 U626 ( .A(n13058), .B(n13018), .C(n359), .Y(n4722) );
  NAND2X1 U627 ( .A(ram[285]), .B(n13018), .Y(n359) );
  OAI21X1 U628 ( .A(n13057), .B(n13018), .C(n360), .Y(n4723) );
  NAND2X1 U629 ( .A(ram[286]), .B(n13018), .Y(n360) );
  OAI21X1 U630 ( .A(n13056), .B(n13018), .C(n361), .Y(n4724) );
  NAND2X1 U631 ( .A(ram[287]), .B(n13018), .Y(n361) );
  OAI21X1 U633 ( .A(n13071), .B(n13017), .C(n363), .Y(n4725) );
  NAND2X1 U634 ( .A(ram[288]), .B(n13017), .Y(n363) );
  OAI21X1 U635 ( .A(n13070), .B(n13017), .C(n364), .Y(n4726) );
  NAND2X1 U636 ( .A(ram[289]), .B(n13017), .Y(n364) );
  OAI21X1 U637 ( .A(n12762), .B(n13017), .C(n365), .Y(n4727) );
  NAND2X1 U638 ( .A(ram[290]), .B(n13017), .Y(n365) );
  OAI21X1 U639 ( .A(n12756), .B(n13017), .C(n366), .Y(n4728) );
  NAND2X1 U640 ( .A(ram[291]), .B(n13017), .Y(n366) );
  OAI21X1 U641 ( .A(n12750), .B(n13017), .C(n367), .Y(n4729) );
  NAND2X1 U642 ( .A(ram[292]), .B(n13017), .Y(n367) );
  OAI21X1 U643 ( .A(n12744), .B(n13017), .C(n368), .Y(n4730) );
  NAND2X1 U644 ( .A(ram[293]), .B(n13017), .Y(n368) );
  OAI21X1 U645 ( .A(n12738), .B(n13017), .C(n369), .Y(n4731) );
  NAND2X1 U646 ( .A(ram[294]), .B(n13017), .Y(n369) );
  OAI21X1 U647 ( .A(n12732), .B(n13017), .C(n370), .Y(n4732) );
  NAND2X1 U648 ( .A(ram[295]), .B(n13017), .Y(n370) );
  OAI21X1 U649 ( .A(n12726), .B(n13017), .C(n371), .Y(n4733) );
  NAND2X1 U650 ( .A(ram[296]), .B(n13017), .Y(n371) );
  OAI21X1 U651 ( .A(n12720), .B(n13017), .C(n372), .Y(n4734) );
  NAND2X1 U652 ( .A(ram[297]), .B(n13017), .Y(n372) );
  OAI21X1 U653 ( .A(n12714), .B(n13017), .C(n373), .Y(n4735) );
  NAND2X1 U654 ( .A(ram[298]), .B(n13017), .Y(n373) );
  OAI21X1 U655 ( .A(n12708), .B(n13017), .C(n374), .Y(n4736) );
  NAND2X1 U656 ( .A(ram[299]), .B(n13017), .Y(n374) );
  OAI21X1 U657 ( .A(n12702), .B(n13017), .C(n375), .Y(n4737) );
  NAND2X1 U658 ( .A(ram[300]), .B(n13017), .Y(n375) );
  OAI21X1 U659 ( .A(n12696), .B(n13017), .C(n376), .Y(n4738) );
  NAND2X1 U660 ( .A(ram[301]), .B(n13017), .Y(n376) );
  OAI21X1 U661 ( .A(n13057), .B(n13017), .C(n377), .Y(n4739) );
  NAND2X1 U662 ( .A(ram[302]), .B(n13017), .Y(n377) );
  OAI21X1 U663 ( .A(n13056), .B(n13017), .C(n378), .Y(n4740) );
  NAND2X1 U664 ( .A(ram[303]), .B(n13017), .Y(n378) );
  OAI21X1 U666 ( .A(n12774), .B(n13016), .C(n380), .Y(n4741) );
  NAND2X1 U667 ( .A(ram[304]), .B(n13016), .Y(n380) );
  OAI21X1 U668 ( .A(n12768), .B(n13016), .C(n381), .Y(n4742) );
  NAND2X1 U669 ( .A(ram[305]), .B(n13016), .Y(n381) );
  OAI21X1 U670 ( .A(n12766), .B(n13016), .C(n382), .Y(n4743) );
  NAND2X1 U671 ( .A(ram[306]), .B(n13016), .Y(n382) );
  OAI21X1 U672 ( .A(n12760), .B(n13016), .C(n383), .Y(n4744) );
  NAND2X1 U673 ( .A(ram[307]), .B(n13016), .Y(n383) );
  OAI21X1 U674 ( .A(n12754), .B(n13016), .C(n384), .Y(n4745) );
  NAND2X1 U675 ( .A(ram[308]), .B(n13016), .Y(n384) );
  OAI21X1 U676 ( .A(n12748), .B(n13016), .C(n385), .Y(n4746) );
  NAND2X1 U677 ( .A(ram[309]), .B(n13016), .Y(n385) );
  OAI21X1 U678 ( .A(n12742), .B(n13016), .C(n386), .Y(n4747) );
  NAND2X1 U679 ( .A(ram[310]), .B(n13016), .Y(n386) );
  OAI21X1 U680 ( .A(n12736), .B(n13016), .C(n387), .Y(n4748) );
  NAND2X1 U681 ( .A(ram[311]), .B(n13016), .Y(n387) );
  OAI21X1 U682 ( .A(n12730), .B(n13016), .C(n388), .Y(n4749) );
  NAND2X1 U683 ( .A(ram[312]), .B(n13016), .Y(n388) );
  OAI21X1 U684 ( .A(n12724), .B(n13016), .C(n389), .Y(n4750) );
  NAND2X1 U685 ( .A(ram[313]), .B(n13016), .Y(n389) );
  OAI21X1 U686 ( .A(n12718), .B(n13016), .C(n390), .Y(n4751) );
  NAND2X1 U687 ( .A(ram[314]), .B(n13016), .Y(n390) );
  OAI21X1 U688 ( .A(n12712), .B(n13016), .C(n391), .Y(n4752) );
  NAND2X1 U689 ( .A(ram[315]), .B(n13016), .Y(n391) );
  OAI21X1 U690 ( .A(n12706), .B(n13016), .C(n392), .Y(n4753) );
  NAND2X1 U691 ( .A(ram[316]), .B(n13016), .Y(n392) );
  OAI21X1 U692 ( .A(n12700), .B(n13016), .C(n393), .Y(n4754) );
  NAND2X1 U693 ( .A(ram[317]), .B(n13016), .Y(n393) );
  OAI21X1 U694 ( .A(n12690), .B(n13016), .C(n394), .Y(n4755) );
  NAND2X1 U695 ( .A(ram[318]), .B(n13016), .Y(n394) );
  OAI21X1 U696 ( .A(n12684), .B(n13016), .C(n395), .Y(n4756) );
  NAND2X1 U697 ( .A(ram[319]), .B(n13016), .Y(n395) );
  OAI21X1 U699 ( .A(n12779), .B(n13015), .C(n397), .Y(n4757) );
  NAND2X1 U700 ( .A(ram[320]), .B(n13015), .Y(n397) );
  OAI21X1 U701 ( .A(n12773), .B(n13015), .C(n398), .Y(n4758) );
  NAND2X1 U702 ( .A(ram[321]), .B(n13015), .Y(n398) );
  OAI21X1 U703 ( .A(n12763), .B(n13015), .C(n399), .Y(n4759) );
  NAND2X1 U704 ( .A(ram[322]), .B(n13015), .Y(n399) );
  OAI21X1 U705 ( .A(n12757), .B(n13015), .C(n400), .Y(n4760) );
  NAND2X1 U706 ( .A(ram[323]), .B(n13015), .Y(n400) );
  OAI21X1 U707 ( .A(n12751), .B(n13015), .C(n401), .Y(n4761) );
  NAND2X1 U708 ( .A(ram[324]), .B(n13015), .Y(n401) );
  OAI21X1 U709 ( .A(n12745), .B(n13015), .C(n402), .Y(n4762) );
  NAND2X1 U710 ( .A(ram[325]), .B(n13015), .Y(n402) );
  OAI21X1 U711 ( .A(n12739), .B(n13015), .C(n403), .Y(n4763) );
  NAND2X1 U712 ( .A(ram[326]), .B(n13015), .Y(n403) );
  OAI21X1 U713 ( .A(n12733), .B(n13015), .C(n404), .Y(n4764) );
  NAND2X1 U714 ( .A(ram[327]), .B(n13015), .Y(n404) );
  OAI21X1 U715 ( .A(n12727), .B(n13015), .C(n405), .Y(n4765) );
  NAND2X1 U716 ( .A(ram[328]), .B(n13015), .Y(n405) );
  OAI21X1 U717 ( .A(n12721), .B(n13015), .C(n406), .Y(n4766) );
  NAND2X1 U718 ( .A(ram[329]), .B(n13015), .Y(n406) );
  OAI21X1 U719 ( .A(n12715), .B(n13015), .C(n407), .Y(n4767) );
  NAND2X1 U720 ( .A(ram[330]), .B(n13015), .Y(n407) );
  OAI21X1 U721 ( .A(n12709), .B(n13015), .C(n408), .Y(n4768) );
  NAND2X1 U722 ( .A(ram[331]), .B(n13015), .Y(n408) );
  OAI21X1 U723 ( .A(n12703), .B(n13015), .C(n409), .Y(n4769) );
  NAND2X1 U724 ( .A(ram[332]), .B(n13015), .Y(n409) );
  OAI21X1 U725 ( .A(n12697), .B(n13015), .C(n410), .Y(n4770) );
  NAND2X1 U726 ( .A(ram[333]), .B(n13015), .Y(n410) );
  OAI21X1 U727 ( .A(n12695), .B(n13015), .C(n411), .Y(n4771) );
  NAND2X1 U728 ( .A(ram[334]), .B(n13015), .Y(n411) );
  OAI21X1 U729 ( .A(n12689), .B(n13015), .C(n412), .Y(n4772) );
  NAND2X1 U730 ( .A(ram[335]), .B(n13015), .Y(n412) );
  OAI21X1 U732 ( .A(n12775), .B(n13014), .C(n414), .Y(n4773) );
  NAND2X1 U733 ( .A(ram[336]), .B(n13014), .Y(n414) );
  OAI21X1 U734 ( .A(n12769), .B(n13014), .C(n415), .Y(n4774) );
  NAND2X1 U735 ( .A(ram[337]), .B(n13014), .Y(n415) );
  OAI21X1 U736 ( .A(n12762), .B(n13014), .C(n416), .Y(n4775) );
  NAND2X1 U737 ( .A(ram[338]), .B(n13014), .Y(n416) );
  OAI21X1 U738 ( .A(n12756), .B(n13014), .C(n417), .Y(n4776) );
  NAND2X1 U739 ( .A(ram[339]), .B(n13014), .Y(n417) );
  OAI21X1 U740 ( .A(n12750), .B(n13014), .C(n418), .Y(n4777) );
  NAND2X1 U741 ( .A(ram[340]), .B(n13014), .Y(n418) );
  OAI21X1 U742 ( .A(n12744), .B(n13014), .C(n419), .Y(n4778) );
  NAND2X1 U743 ( .A(ram[341]), .B(n13014), .Y(n419) );
  OAI21X1 U744 ( .A(n12738), .B(n13014), .C(n420), .Y(n4779) );
  NAND2X1 U745 ( .A(ram[342]), .B(n13014), .Y(n420) );
  OAI21X1 U746 ( .A(n12732), .B(n13014), .C(n421), .Y(n4780) );
  NAND2X1 U747 ( .A(ram[343]), .B(n13014), .Y(n421) );
  OAI21X1 U748 ( .A(n12726), .B(n13014), .C(n422), .Y(n4781) );
  NAND2X1 U749 ( .A(ram[344]), .B(n13014), .Y(n422) );
  OAI21X1 U750 ( .A(n12720), .B(n13014), .C(n423), .Y(n4782) );
  NAND2X1 U751 ( .A(ram[345]), .B(n13014), .Y(n423) );
  OAI21X1 U752 ( .A(n12714), .B(n13014), .C(n424), .Y(n4783) );
  NAND2X1 U753 ( .A(ram[346]), .B(n13014), .Y(n424) );
  OAI21X1 U754 ( .A(n12708), .B(n13014), .C(n425), .Y(n4784) );
  NAND2X1 U755 ( .A(ram[347]), .B(n13014), .Y(n425) );
  OAI21X1 U756 ( .A(n12702), .B(n13014), .C(n426), .Y(n4785) );
  NAND2X1 U757 ( .A(ram[348]), .B(n13014), .Y(n426) );
  OAI21X1 U758 ( .A(n12696), .B(n13014), .C(n427), .Y(n4786) );
  NAND2X1 U759 ( .A(ram[349]), .B(n13014), .Y(n427) );
  OAI21X1 U760 ( .A(n12691), .B(n13014), .C(n428), .Y(n4787) );
  NAND2X1 U761 ( .A(ram[350]), .B(n13014), .Y(n428) );
  OAI21X1 U762 ( .A(n12685), .B(n13014), .C(n429), .Y(n4788) );
  NAND2X1 U763 ( .A(ram[351]), .B(n13014), .Y(n429) );
  OAI21X1 U765 ( .A(n12778), .B(n13013), .C(n431), .Y(n4789) );
  NAND2X1 U766 ( .A(ram[352]), .B(n13013), .Y(n431) );
  OAI21X1 U767 ( .A(n12772), .B(n13013), .C(n432), .Y(n4790) );
  NAND2X1 U768 ( .A(ram[353]), .B(n13013), .Y(n432) );
  OAI21X1 U769 ( .A(n12762), .B(n13013), .C(n433), .Y(n4791) );
  NAND2X1 U770 ( .A(ram[354]), .B(n13013), .Y(n433) );
  OAI21X1 U771 ( .A(n12756), .B(n13013), .C(n434), .Y(n4792) );
  NAND2X1 U772 ( .A(ram[355]), .B(n13013), .Y(n434) );
  OAI21X1 U773 ( .A(n12750), .B(n13013), .C(n435), .Y(n4793) );
  NAND2X1 U774 ( .A(ram[356]), .B(n13013), .Y(n435) );
  OAI21X1 U775 ( .A(n12744), .B(n13013), .C(n436), .Y(n4794) );
  NAND2X1 U776 ( .A(ram[357]), .B(n13013), .Y(n436) );
  OAI21X1 U777 ( .A(n12738), .B(n13013), .C(n437), .Y(n4795) );
  NAND2X1 U778 ( .A(ram[358]), .B(n13013), .Y(n437) );
  OAI21X1 U779 ( .A(n12732), .B(n13013), .C(n438), .Y(n4796) );
  NAND2X1 U780 ( .A(ram[359]), .B(n13013), .Y(n438) );
  OAI21X1 U781 ( .A(n12726), .B(n13013), .C(n439), .Y(n4797) );
  NAND2X1 U782 ( .A(ram[360]), .B(n13013), .Y(n439) );
  OAI21X1 U783 ( .A(n12720), .B(n13013), .C(n440), .Y(n4798) );
  NAND2X1 U784 ( .A(ram[361]), .B(n13013), .Y(n440) );
  OAI21X1 U785 ( .A(n12714), .B(n13013), .C(n441), .Y(n4799) );
  NAND2X1 U786 ( .A(ram[362]), .B(n13013), .Y(n441) );
  OAI21X1 U787 ( .A(n12708), .B(n13013), .C(n442), .Y(n4800) );
  NAND2X1 U788 ( .A(ram[363]), .B(n13013), .Y(n442) );
  OAI21X1 U789 ( .A(n12702), .B(n13013), .C(n443), .Y(n4801) );
  NAND2X1 U790 ( .A(ram[364]), .B(n13013), .Y(n443) );
  OAI21X1 U791 ( .A(n12696), .B(n13013), .C(n444), .Y(n4802) );
  NAND2X1 U792 ( .A(ram[365]), .B(n13013), .Y(n444) );
  OAI21X1 U793 ( .A(n12694), .B(n13013), .C(n445), .Y(n4803) );
  NAND2X1 U794 ( .A(ram[366]), .B(n13013), .Y(n445) );
  OAI21X1 U795 ( .A(n12688), .B(n13013), .C(n446), .Y(n4804) );
  NAND2X1 U796 ( .A(ram[367]), .B(n13013), .Y(n446) );
  OAI21X1 U798 ( .A(n12779), .B(n13012), .C(n448), .Y(n4805) );
  NAND2X1 U799 ( .A(ram[368]), .B(n13012), .Y(n448) );
  OAI21X1 U800 ( .A(n12773), .B(n13012), .C(n449), .Y(n4806) );
  NAND2X1 U801 ( .A(ram[369]), .B(n13012), .Y(n449) );
  OAI21X1 U802 ( .A(n12763), .B(n13012), .C(n450), .Y(n4807) );
  NAND2X1 U803 ( .A(ram[370]), .B(n13012), .Y(n450) );
  OAI21X1 U804 ( .A(n12757), .B(n13012), .C(n451), .Y(n4808) );
  NAND2X1 U805 ( .A(ram[371]), .B(n13012), .Y(n451) );
  OAI21X1 U806 ( .A(n12751), .B(n13012), .C(n452), .Y(n4809) );
  NAND2X1 U807 ( .A(ram[372]), .B(n13012), .Y(n452) );
  OAI21X1 U808 ( .A(n12745), .B(n13012), .C(n453), .Y(n4810) );
  NAND2X1 U809 ( .A(ram[373]), .B(n13012), .Y(n453) );
  OAI21X1 U810 ( .A(n12739), .B(n13012), .C(n454), .Y(n4811) );
  NAND2X1 U811 ( .A(ram[374]), .B(n13012), .Y(n454) );
  OAI21X1 U812 ( .A(n12733), .B(n13012), .C(n455), .Y(n4812) );
  NAND2X1 U813 ( .A(ram[375]), .B(n13012), .Y(n455) );
  OAI21X1 U814 ( .A(n12727), .B(n13012), .C(n456), .Y(n4813) );
  NAND2X1 U815 ( .A(ram[376]), .B(n13012), .Y(n456) );
  OAI21X1 U816 ( .A(n12721), .B(n13012), .C(n457), .Y(n4814) );
  NAND2X1 U817 ( .A(ram[377]), .B(n13012), .Y(n457) );
  OAI21X1 U818 ( .A(n12715), .B(n13012), .C(n458), .Y(n4815) );
  NAND2X1 U819 ( .A(ram[378]), .B(n13012), .Y(n458) );
  OAI21X1 U820 ( .A(n12709), .B(n13012), .C(n459), .Y(n4816) );
  NAND2X1 U821 ( .A(ram[379]), .B(n13012), .Y(n459) );
  OAI21X1 U822 ( .A(n12703), .B(n13012), .C(n460), .Y(n4817) );
  NAND2X1 U823 ( .A(ram[380]), .B(n13012), .Y(n460) );
  OAI21X1 U824 ( .A(n12697), .B(n13012), .C(n461), .Y(n4818) );
  NAND2X1 U825 ( .A(ram[381]), .B(n13012), .Y(n461) );
  OAI21X1 U826 ( .A(n12695), .B(n13012), .C(n462), .Y(n4819) );
  NAND2X1 U827 ( .A(ram[382]), .B(n13012), .Y(n462) );
  OAI21X1 U828 ( .A(n12689), .B(n13012), .C(n463), .Y(n4820) );
  NAND2X1 U829 ( .A(ram[383]), .B(n13012), .Y(n463) );
  OAI21X1 U831 ( .A(n12774), .B(n13011), .C(n465), .Y(n4821) );
  NAND2X1 U832 ( .A(ram[384]), .B(n13011), .Y(n465) );
  OAI21X1 U833 ( .A(n12768), .B(n13011), .C(n466), .Y(n4822) );
  NAND2X1 U834 ( .A(ram[385]), .B(n13011), .Y(n466) );
  OAI21X1 U835 ( .A(n12763), .B(n13011), .C(n467), .Y(n4823) );
  NAND2X1 U836 ( .A(ram[386]), .B(n13011), .Y(n467) );
  OAI21X1 U837 ( .A(n12757), .B(n13011), .C(n468), .Y(n4824) );
  NAND2X1 U838 ( .A(ram[387]), .B(n13011), .Y(n468) );
  OAI21X1 U839 ( .A(n12751), .B(n13011), .C(n469), .Y(n4825) );
  NAND2X1 U840 ( .A(ram[388]), .B(n13011), .Y(n469) );
  OAI21X1 U841 ( .A(n12745), .B(n13011), .C(n470), .Y(n4826) );
  NAND2X1 U842 ( .A(ram[389]), .B(n13011), .Y(n470) );
  OAI21X1 U843 ( .A(n12739), .B(n13011), .C(n471), .Y(n4827) );
  NAND2X1 U844 ( .A(ram[390]), .B(n13011), .Y(n471) );
  OAI21X1 U845 ( .A(n12733), .B(n13011), .C(n472), .Y(n4828) );
  NAND2X1 U846 ( .A(ram[391]), .B(n13011), .Y(n472) );
  OAI21X1 U847 ( .A(n12727), .B(n13011), .C(n473), .Y(n4829) );
  NAND2X1 U848 ( .A(ram[392]), .B(n13011), .Y(n473) );
  OAI21X1 U849 ( .A(n12721), .B(n13011), .C(n474), .Y(n4830) );
  NAND2X1 U850 ( .A(ram[393]), .B(n13011), .Y(n474) );
  OAI21X1 U851 ( .A(n12715), .B(n13011), .C(n475), .Y(n4831) );
  NAND2X1 U852 ( .A(ram[394]), .B(n13011), .Y(n475) );
  OAI21X1 U853 ( .A(n12709), .B(n13011), .C(n476), .Y(n4832) );
  NAND2X1 U854 ( .A(ram[395]), .B(n13011), .Y(n476) );
  OAI21X1 U855 ( .A(n12703), .B(n13011), .C(n477), .Y(n4833) );
  NAND2X1 U856 ( .A(ram[396]), .B(n13011), .Y(n477) );
  OAI21X1 U857 ( .A(n12697), .B(n13011), .C(n478), .Y(n4834) );
  NAND2X1 U858 ( .A(ram[397]), .B(n13011), .Y(n478) );
  OAI21X1 U859 ( .A(n12690), .B(n13011), .C(n479), .Y(n4835) );
  NAND2X1 U860 ( .A(ram[398]), .B(n13011), .Y(n479) );
  OAI21X1 U861 ( .A(n12684), .B(n13011), .C(n480), .Y(n4836) );
  NAND2X1 U862 ( .A(ram[399]), .B(n13011), .Y(n480) );
  OAI21X1 U864 ( .A(n12775), .B(n13010), .C(n482), .Y(n4837) );
  NAND2X1 U865 ( .A(ram[400]), .B(n13010), .Y(n482) );
  OAI21X1 U866 ( .A(n12769), .B(n13010), .C(n483), .Y(n4838) );
  NAND2X1 U867 ( .A(ram[401]), .B(n13010), .Y(n483) );
  OAI21X1 U868 ( .A(n12765), .B(n13010), .C(n484), .Y(n4839) );
  NAND2X1 U869 ( .A(ram[402]), .B(n13010), .Y(n484) );
  OAI21X1 U870 ( .A(n12759), .B(n13010), .C(n485), .Y(n4840) );
  NAND2X1 U871 ( .A(ram[403]), .B(n13010), .Y(n485) );
  OAI21X1 U872 ( .A(n12753), .B(n13010), .C(n486), .Y(n4841) );
  NAND2X1 U873 ( .A(ram[404]), .B(n13010), .Y(n486) );
  OAI21X1 U874 ( .A(n12747), .B(n13010), .C(n487), .Y(n4842) );
  NAND2X1 U875 ( .A(ram[405]), .B(n13010), .Y(n487) );
  OAI21X1 U876 ( .A(n12741), .B(n13010), .C(n488), .Y(n4843) );
  NAND2X1 U877 ( .A(ram[406]), .B(n13010), .Y(n488) );
  OAI21X1 U878 ( .A(n12735), .B(n13010), .C(n489), .Y(n4844) );
  NAND2X1 U879 ( .A(ram[407]), .B(n13010), .Y(n489) );
  OAI21X1 U880 ( .A(n12729), .B(n13010), .C(n490), .Y(n4845) );
  NAND2X1 U881 ( .A(ram[408]), .B(n13010), .Y(n490) );
  OAI21X1 U882 ( .A(n12723), .B(n13010), .C(n491), .Y(n4846) );
  NAND2X1 U883 ( .A(ram[409]), .B(n13010), .Y(n491) );
  OAI21X1 U884 ( .A(n12717), .B(n13010), .C(n492), .Y(n4847) );
  NAND2X1 U885 ( .A(ram[410]), .B(n13010), .Y(n492) );
  OAI21X1 U886 ( .A(n12711), .B(n13010), .C(n493), .Y(n4848) );
  NAND2X1 U887 ( .A(ram[411]), .B(n13010), .Y(n493) );
  OAI21X1 U888 ( .A(n12705), .B(n13010), .C(n494), .Y(n4849) );
  NAND2X1 U889 ( .A(ram[412]), .B(n13010), .Y(n494) );
  OAI21X1 U890 ( .A(n12699), .B(n13010), .C(n495), .Y(n4850) );
  NAND2X1 U891 ( .A(ram[413]), .B(n13010), .Y(n495) );
  OAI21X1 U892 ( .A(n12691), .B(n13010), .C(n496), .Y(n4851) );
  NAND2X1 U893 ( .A(ram[414]), .B(n13010), .Y(n496) );
  OAI21X1 U894 ( .A(n12685), .B(n13010), .C(n497), .Y(n4852) );
  NAND2X1 U895 ( .A(ram[415]), .B(n13010), .Y(n497) );
  OAI21X1 U897 ( .A(n12774), .B(n13009), .C(n499), .Y(n4853) );
  NAND2X1 U898 ( .A(ram[416]), .B(n13009), .Y(n499) );
  OAI21X1 U899 ( .A(n12768), .B(n13009), .C(n500), .Y(n4854) );
  NAND2X1 U900 ( .A(ram[417]), .B(n13009), .Y(n500) );
  OAI21X1 U901 ( .A(n12762), .B(n13009), .C(n501), .Y(n4855) );
  NAND2X1 U902 ( .A(ram[418]), .B(n13009), .Y(n501) );
  OAI21X1 U903 ( .A(n12756), .B(n13009), .C(n502), .Y(n4856) );
  NAND2X1 U904 ( .A(ram[419]), .B(n13009), .Y(n502) );
  OAI21X1 U905 ( .A(n12750), .B(n13009), .C(n503), .Y(n4857) );
  NAND2X1 U906 ( .A(ram[420]), .B(n13009), .Y(n503) );
  OAI21X1 U907 ( .A(n12744), .B(n13009), .C(n504), .Y(n4858) );
  NAND2X1 U908 ( .A(ram[421]), .B(n13009), .Y(n504) );
  OAI21X1 U909 ( .A(n12738), .B(n13009), .C(n505), .Y(n4859) );
  NAND2X1 U910 ( .A(ram[422]), .B(n13009), .Y(n505) );
  OAI21X1 U911 ( .A(n12732), .B(n13009), .C(n506), .Y(n4860) );
  NAND2X1 U912 ( .A(ram[423]), .B(n13009), .Y(n506) );
  OAI21X1 U913 ( .A(n12726), .B(n13009), .C(n507), .Y(n4861) );
  NAND2X1 U914 ( .A(ram[424]), .B(n13009), .Y(n507) );
  OAI21X1 U915 ( .A(n12720), .B(n13009), .C(n508), .Y(n4862) );
  NAND2X1 U916 ( .A(ram[425]), .B(n13009), .Y(n508) );
  OAI21X1 U917 ( .A(n12714), .B(n13009), .C(n509), .Y(n4863) );
  NAND2X1 U918 ( .A(ram[426]), .B(n13009), .Y(n509) );
  OAI21X1 U919 ( .A(n12708), .B(n13009), .C(n510), .Y(n4864) );
  NAND2X1 U920 ( .A(ram[427]), .B(n13009), .Y(n510) );
  OAI21X1 U921 ( .A(n12702), .B(n13009), .C(n511), .Y(n4865) );
  NAND2X1 U922 ( .A(ram[428]), .B(n13009), .Y(n511) );
  OAI21X1 U923 ( .A(n12696), .B(n13009), .C(n512), .Y(n4866) );
  NAND2X1 U924 ( .A(ram[429]), .B(n13009), .Y(n512) );
  OAI21X1 U925 ( .A(n12690), .B(n13009), .C(n513), .Y(n4867) );
  NAND2X1 U926 ( .A(ram[430]), .B(n13009), .Y(n513) );
  OAI21X1 U927 ( .A(n12684), .B(n13009), .C(n514), .Y(n4868) );
  NAND2X1 U928 ( .A(ram[431]), .B(n13009), .Y(n514) );
  OAI21X1 U930 ( .A(n12774), .B(n13008), .C(n516), .Y(n4869) );
  NAND2X1 U931 ( .A(ram[432]), .B(n13008), .Y(n516) );
  OAI21X1 U932 ( .A(n12768), .B(n13008), .C(n517), .Y(n4870) );
  NAND2X1 U933 ( .A(ram[433]), .B(n13008), .Y(n517) );
  OAI21X1 U934 ( .A(n12767), .B(n13008), .C(n518), .Y(n4871) );
  NAND2X1 U935 ( .A(ram[434]), .B(n13008), .Y(n518) );
  OAI21X1 U936 ( .A(n12761), .B(n13008), .C(n519), .Y(n4872) );
  NAND2X1 U937 ( .A(ram[435]), .B(n13008), .Y(n519) );
  OAI21X1 U938 ( .A(n12755), .B(n13008), .C(n520), .Y(n4873) );
  NAND2X1 U939 ( .A(ram[436]), .B(n13008), .Y(n520) );
  OAI21X1 U940 ( .A(n12749), .B(n13008), .C(n521), .Y(n4874) );
  NAND2X1 U941 ( .A(ram[437]), .B(n13008), .Y(n521) );
  OAI21X1 U942 ( .A(n12743), .B(n13008), .C(n522), .Y(n4875) );
  NAND2X1 U943 ( .A(ram[438]), .B(n13008), .Y(n522) );
  OAI21X1 U944 ( .A(n12737), .B(n13008), .C(n523), .Y(n4876) );
  NAND2X1 U945 ( .A(ram[439]), .B(n13008), .Y(n523) );
  OAI21X1 U946 ( .A(n12731), .B(n13008), .C(n524), .Y(n4877) );
  NAND2X1 U947 ( .A(ram[440]), .B(n13008), .Y(n524) );
  OAI21X1 U948 ( .A(n12725), .B(n13008), .C(n525), .Y(n4878) );
  NAND2X1 U949 ( .A(ram[441]), .B(n13008), .Y(n525) );
  OAI21X1 U950 ( .A(n12719), .B(n13008), .C(n526), .Y(n4879) );
  NAND2X1 U951 ( .A(ram[442]), .B(n13008), .Y(n526) );
  OAI21X1 U952 ( .A(n12713), .B(n13008), .C(n527), .Y(n4880) );
  NAND2X1 U953 ( .A(ram[443]), .B(n13008), .Y(n527) );
  OAI21X1 U954 ( .A(n12707), .B(n13008), .C(n528), .Y(n4881) );
  NAND2X1 U955 ( .A(ram[444]), .B(n13008), .Y(n528) );
  OAI21X1 U956 ( .A(n12701), .B(n13008), .C(n529), .Y(n4882) );
  NAND2X1 U957 ( .A(ram[445]), .B(n13008), .Y(n529) );
  OAI21X1 U958 ( .A(n12690), .B(n13008), .C(n530), .Y(n4883) );
  NAND2X1 U959 ( .A(ram[446]), .B(n13008), .Y(n530) );
  OAI21X1 U960 ( .A(n12684), .B(n13008), .C(n531), .Y(n4884) );
  NAND2X1 U961 ( .A(ram[447]), .B(n13008), .Y(n531) );
  OAI21X1 U963 ( .A(n12775), .B(n13007), .C(n533), .Y(n4885) );
  NAND2X1 U964 ( .A(ram[448]), .B(n13007), .Y(n533) );
  OAI21X1 U965 ( .A(n12769), .B(n13007), .C(n534), .Y(n4886) );
  NAND2X1 U966 ( .A(ram[449]), .B(n13007), .Y(n534) );
  OAI21X1 U967 ( .A(n12762), .B(n13007), .C(n535), .Y(n4887) );
  NAND2X1 U968 ( .A(ram[450]), .B(n13007), .Y(n535) );
  OAI21X1 U969 ( .A(n12756), .B(n13007), .C(n536), .Y(n4888) );
  NAND2X1 U970 ( .A(ram[451]), .B(n13007), .Y(n536) );
  OAI21X1 U971 ( .A(n12750), .B(n13007), .C(n537), .Y(n4889) );
  NAND2X1 U972 ( .A(ram[452]), .B(n13007), .Y(n537) );
  OAI21X1 U973 ( .A(n12744), .B(n13007), .C(n538), .Y(n4890) );
  NAND2X1 U974 ( .A(ram[453]), .B(n13007), .Y(n538) );
  OAI21X1 U975 ( .A(n12738), .B(n13007), .C(n539), .Y(n4891) );
  NAND2X1 U976 ( .A(ram[454]), .B(n13007), .Y(n539) );
  OAI21X1 U977 ( .A(n12732), .B(n13007), .C(n540), .Y(n4892) );
  NAND2X1 U978 ( .A(ram[455]), .B(n13007), .Y(n540) );
  OAI21X1 U979 ( .A(n12726), .B(n13007), .C(n541), .Y(n4893) );
  NAND2X1 U980 ( .A(ram[456]), .B(n13007), .Y(n541) );
  OAI21X1 U981 ( .A(n12720), .B(n13007), .C(n542), .Y(n4894) );
  NAND2X1 U982 ( .A(ram[457]), .B(n13007), .Y(n542) );
  OAI21X1 U983 ( .A(n12714), .B(n13007), .C(n543), .Y(n4895) );
  NAND2X1 U984 ( .A(ram[458]), .B(n13007), .Y(n543) );
  OAI21X1 U985 ( .A(n12708), .B(n13007), .C(n544), .Y(n4896) );
  NAND2X1 U986 ( .A(ram[459]), .B(n13007), .Y(n544) );
  OAI21X1 U987 ( .A(n12702), .B(n13007), .C(n545), .Y(n4897) );
  NAND2X1 U988 ( .A(ram[460]), .B(n13007), .Y(n545) );
  OAI21X1 U989 ( .A(n12696), .B(n13007), .C(n546), .Y(n4898) );
  NAND2X1 U990 ( .A(ram[461]), .B(n13007), .Y(n546) );
  OAI21X1 U991 ( .A(n12691), .B(n13007), .C(n547), .Y(n4899) );
  NAND2X1 U992 ( .A(ram[462]), .B(n13007), .Y(n547) );
  OAI21X1 U993 ( .A(n12685), .B(n13007), .C(n548), .Y(n4900) );
  NAND2X1 U994 ( .A(ram[463]), .B(n13007), .Y(n548) );
  OAI21X1 U996 ( .A(n12774), .B(n13006), .C(n550), .Y(n4901) );
  NAND2X1 U997 ( .A(ram[464]), .B(n13006), .Y(n550) );
  OAI21X1 U998 ( .A(n12768), .B(n13006), .C(n551), .Y(n4902) );
  NAND2X1 U999 ( .A(ram[465]), .B(n13006), .Y(n551) );
  OAI21X1 U1000 ( .A(n12764), .B(n13006), .C(n552), .Y(n4903) );
  NAND2X1 U1001 ( .A(ram[466]), .B(n13006), .Y(n552) );
  OAI21X1 U1002 ( .A(n12758), .B(n13006), .C(n553), .Y(n4904) );
  NAND2X1 U1003 ( .A(ram[467]), .B(n13006), .Y(n553) );
  OAI21X1 U1004 ( .A(n12752), .B(n13006), .C(n554), .Y(n4905) );
  NAND2X1 U1005 ( .A(ram[468]), .B(n13006), .Y(n554) );
  OAI21X1 U1006 ( .A(n12746), .B(n13006), .C(n555), .Y(n4906) );
  NAND2X1 U1007 ( .A(ram[469]), .B(n13006), .Y(n555) );
  OAI21X1 U1008 ( .A(n12740), .B(n13006), .C(n556), .Y(n4907) );
  NAND2X1 U1009 ( .A(ram[470]), .B(n13006), .Y(n556) );
  OAI21X1 U1010 ( .A(n12734), .B(n13006), .C(n557), .Y(n4908) );
  NAND2X1 U1011 ( .A(ram[471]), .B(n13006), .Y(n557) );
  OAI21X1 U1012 ( .A(n12728), .B(n13006), .C(n558), .Y(n4909) );
  NAND2X1 U1013 ( .A(ram[472]), .B(n13006), .Y(n558) );
  OAI21X1 U1014 ( .A(n12722), .B(n13006), .C(n559), .Y(n4910) );
  NAND2X1 U1015 ( .A(ram[473]), .B(n13006), .Y(n559) );
  OAI21X1 U1016 ( .A(n12716), .B(n13006), .C(n560), .Y(n4911) );
  NAND2X1 U1017 ( .A(ram[474]), .B(n13006), .Y(n560) );
  OAI21X1 U1018 ( .A(n12710), .B(n13006), .C(n561), .Y(n4912) );
  NAND2X1 U1019 ( .A(ram[475]), .B(n13006), .Y(n561) );
  OAI21X1 U1020 ( .A(n12704), .B(n13006), .C(n562), .Y(n4913) );
  NAND2X1 U1021 ( .A(ram[476]), .B(n13006), .Y(n562) );
  OAI21X1 U1022 ( .A(n12698), .B(n13006), .C(n563), .Y(n4914) );
  NAND2X1 U1023 ( .A(ram[477]), .B(n13006), .Y(n563) );
  OAI21X1 U1024 ( .A(n12690), .B(n13006), .C(n564), .Y(n4915) );
  NAND2X1 U1025 ( .A(ram[478]), .B(n13006), .Y(n564) );
  OAI21X1 U1026 ( .A(n12684), .B(n13006), .C(n565), .Y(n4916) );
  NAND2X1 U1027 ( .A(ram[479]), .B(n13006), .Y(n565) );
  OAI21X1 U1029 ( .A(n12774), .B(n13005), .C(n567), .Y(n4917) );
  NAND2X1 U1030 ( .A(ram[480]), .B(n13005), .Y(n567) );
  OAI21X1 U1031 ( .A(n12768), .B(n13005), .C(n568), .Y(n4918) );
  NAND2X1 U1032 ( .A(ram[481]), .B(n13005), .Y(n568) );
  OAI21X1 U1033 ( .A(n12762), .B(n13005), .C(n569), .Y(n4919) );
  NAND2X1 U1034 ( .A(ram[482]), .B(n13005), .Y(n569) );
  OAI21X1 U1035 ( .A(n12756), .B(n13005), .C(n570), .Y(n4920) );
  NAND2X1 U1036 ( .A(ram[483]), .B(n13005), .Y(n570) );
  OAI21X1 U1037 ( .A(n12750), .B(n13005), .C(n571), .Y(n4921) );
  NAND2X1 U1038 ( .A(ram[484]), .B(n13005), .Y(n571) );
  OAI21X1 U1039 ( .A(n12744), .B(n13005), .C(n572), .Y(n4922) );
  NAND2X1 U1040 ( .A(ram[485]), .B(n13005), .Y(n572) );
  OAI21X1 U1041 ( .A(n12738), .B(n13005), .C(n573), .Y(n4923) );
  NAND2X1 U1042 ( .A(ram[486]), .B(n13005), .Y(n573) );
  OAI21X1 U1043 ( .A(n12732), .B(n13005), .C(n574), .Y(n4924) );
  NAND2X1 U1044 ( .A(ram[487]), .B(n13005), .Y(n574) );
  OAI21X1 U1045 ( .A(n12726), .B(n13005), .C(n575), .Y(n4925) );
  NAND2X1 U1046 ( .A(ram[488]), .B(n13005), .Y(n575) );
  OAI21X1 U1047 ( .A(n12720), .B(n13005), .C(n576), .Y(n4926) );
  NAND2X1 U1048 ( .A(ram[489]), .B(n13005), .Y(n576) );
  OAI21X1 U1049 ( .A(n12714), .B(n13005), .C(n577), .Y(n4927) );
  NAND2X1 U1050 ( .A(ram[490]), .B(n13005), .Y(n577) );
  OAI21X1 U1051 ( .A(n12708), .B(n13005), .C(n578), .Y(n4928) );
  NAND2X1 U1052 ( .A(ram[491]), .B(n13005), .Y(n578) );
  OAI21X1 U1053 ( .A(n12702), .B(n13005), .C(n579), .Y(n4929) );
  NAND2X1 U1054 ( .A(ram[492]), .B(n13005), .Y(n579) );
  OAI21X1 U1055 ( .A(n12696), .B(n13005), .C(n580), .Y(n4930) );
  NAND2X1 U1056 ( .A(ram[493]), .B(n13005), .Y(n580) );
  OAI21X1 U1057 ( .A(n12690), .B(n13005), .C(n581), .Y(n4931) );
  NAND2X1 U1058 ( .A(ram[494]), .B(n13005), .Y(n581) );
  OAI21X1 U1059 ( .A(n12684), .B(n13005), .C(n582), .Y(n4932) );
  NAND2X1 U1060 ( .A(ram[495]), .B(n13005), .Y(n582) );
  OAI21X1 U1062 ( .A(n12778), .B(n13004), .C(n584), .Y(n4933) );
  NAND2X1 U1063 ( .A(ram[496]), .B(n13004), .Y(n584) );
  OAI21X1 U1064 ( .A(n12772), .B(n13004), .C(n585), .Y(n4934) );
  NAND2X1 U1065 ( .A(ram[497]), .B(n13004), .Y(n585) );
  OAI21X1 U1066 ( .A(n12763), .B(n13004), .C(n586), .Y(n4935) );
  NAND2X1 U1067 ( .A(ram[498]), .B(n13004), .Y(n586) );
  OAI21X1 U1068 ( .A(n12757), .B(n13004), .C(n587), .Y(n4936) );
  NAND2X1 U1069 ( .A(ram[499]), .B(n13004), .Y(n587) );
  OAI21X1 U1070 ( .A(n12751), .B(n13004), .C(n588), .Y(n4937) );
  NAND2X1 U1071 ( .A(ram[500]), .B(n13004), .Y(n588) );
  OAI21X1 U1072 ( .A(n12745), .B(n13004), .C(n589), .Y(n4938) );
  NAND2X1 U1073 ( .A(ram[501]), .B(n13004), .Y(n589) );
  OAI21X1 U1074 ( .A(n12739), .B(n13004), .C(n590), .Y(n4939) );
  NAND2X1 U1075 ( .A(ram[502]), .B(n13004), .Y(n590) );
  OAI21X1 U1076 ( .A(n12733), .B(n13004), .C(n591), .Y(n4940) );
  NAND2X1 U1077 ( .A(ram[503]), .B(n13004), .Y(n591) );
  OAI21X1 U1078 ( .A(n12727), .B(n13004), .C(n592), .Y(n4941) );
  NAND2X1 U1079 ( .A(ram[504]), .B(n13004), .Y(n592) );
  OAI21X1 U1080 ( .A(n12721), .B(n13004), .C(n593), .Y(n4942) );
  NAND2X1 U1081 ( .A(ram[505]), .B(n13004), .Y(n593) );
  OAI21X1 U1082 ( .A(n12715), .B(n13004), .C(n594), .Y(n4943) );
  NAND2X1 U1083 ( .A(ram[506]), .B(n13004), .Y(n594) );
  OAI21X1 U1084 ( .A(n12709), .B(n13004), .C(n595), .Y(n4944) );
  NAND2X1 U1085 ( .A(ram[507]), .B(n13004), .Y(n595) );
  OAI21X1 U1086 ( .A(n12703), .B(n13004), .C(n596), .Y(n4945) );
  NAND2X1 U1087 ( .A(ram[508]), .B(n13004), .Y(n596) );
  OAI21X1 U1088 ( .A(n12697), .B(n13004), .C(n597), .Y(n4946) );
  NAND2X1 U1089 ( .A(ram[509]), .B(n13004), .Y(n597) );
  OAI21X1 U1090 ( .A(n12694), .B(n13004), .C(n598), .Y(n4947) );
  NAND2X1 U1091 ( .A(ram[510]), .B(n13004), .Y(n598) );
  OAI21X1 U1092 ( .A(n12688), .B(n13004), .C(n599), .Y(n4948) );
  NAND2X1 U1093 ( .A(ram[511]), .B(n13004), .Y(n599) );
  NAND3X1 U1095 ( .A(mem_write_en), .B(n326), .C(n601), .Y(n600) );
  OAI21X1 U1096 ( .A(n12775), .B(n13003), .C(n603), .Y(n4949) );
  NAND2X1 U1097 ( .A(ram[512]), .B(n13003), .Y(n603) );
  OAI21X1 U1098 ( .A(n12769), .B(n13003), .C(n604), .Y(n4950) );
  NAND2X1 U1099 ( .A(ram[513]), .B(n13003), .Y(n604) );
  OAI21X1 U1100 ( .A(n12763), .B(n13003), .C(n605), .Y(n4951) );
  NAND2X1 U1101 ( .A(ram[514]), .B(n13003), .Y(n605) );
  OAI21X1 U1102 ( .A(n12757), .B(n13003), .C(n606), .Y(n4952) );
  NAND2X1 U1103 ( .A(ram[515]), .B(n13003), .Y(n606) );
  OAI21X1 U1104 ( .A(n12751), .B(n13003), .C(n607), .Y(n4953) );
  NAND2X1 U1105 ( .A(ram[516]), .B(n13003), .Y(n607) );
  OAI21X1 U1106 ( .A(n12745), .B(n13003), .C(n608), .Y(n4954) );
  NAND2X1 U1107 ( .A(ram[517]), .B(n13003), .Y(n608) );
  OAI21X1 U1108 ( .A(n12739), .B(n13003), .C(n609), .Y(n4955) );
  NAND2X1 U1109 ( .A(ram[518]), .B(n13003), .Y(n609) );
  OAI21X1 U1110 ( .A(n12733), .B(n13003), .C(n610), .Y(n4956) );
  NAND2X1 U1111 ( .A(ram[519]), .B(n13003), .Y(n610) );
  OAI21X1 U1112 ( .A(n12727), .B(n13003), .C(n611), .Y(n4957) );
  NAND2X1 U1113 ( .A(ram[520]), .B(n13003), .Y(n611) );
  OAI21X1 U1114 ( .A(n12721), .B(n13003), .C(n612), .Y(n4958) );
  NAND2X1 U1115 ( .A(ram[521]), .B(n13003), .Y(n612) );
  OAI21X1 U1116 ( .A(n12715), .B(n13003), .C(n613), .Y(n4959) );
  NAND2X1 U1117 ( .A(ram[522]), .B(n13003), .Y(n613) );
  OAI21X1 U1118 ( .A(n12709), .B(n13003), .C(n614), .Y(n4960) );
  NAND2X1 U1119 ( .A(ram[523]), .B(n13003), .Y(n614) );
  OAI21X1 U1120 ( .A(n12703), .B(n13003), .C(n615), .Y(n4961) );
  NAND2X1 U1121 ( .A(ram[524]), .B(n13003), .Y(n615) );
  OAI21X1 U1122 ( .A(n12697), .B(n13003), .C(n616), .Y(n4962) );
  NAND2X1 U1123 ( .A(ram[525]), .B(n13003), .Y(n616) );
  OAI21X1 U1124 ( .A(n12691), .B(n13003), .C(n617), .Y(n4963) );
  NAND2X1 U1125 ( .A(ram[526]), .B(n13003), .Y(n617) );
  OAI21X1 U1126 ( .A(n12685), .B(n13003), .C(n618), .Y(n4964) );
  NAND2X1 U1127 ( .A(ram[527]), .B(n13003), .Y(n618) );
  OAI21X1 U1129 ( .A(n12774), .B(n13002), .C(n620), .Y(n4965) );
  NAND2X1 U1130 ( .A(ram[528]), .B(n13002), .Y(n620) );
  OAI21X1 U1131 ( .A(n12768), .B(n13002), .C(n621), .Y(n4966) );
  NAND2X1 U1132 ( .A(ram[529]), .B(n13002), .Y(n621) );
  OAI21X1 U1133 ( .A(n12762), .B(n13002), .C(n622), .Y(n4967) );
  NAND2X1 U1134 ( .A(ram[530]), .B(n13002), .Y(n622) );
  OAI21X1 U1135 ( .A(n12756), .B(n13002), .C(n623), .Y(n4968) );
  NAND2X1 U1136 ( .A(ram[531]), .B(n13002), .Y(n623) );
  OAI21X1 U1137 ( .A(n12750), .B(n13002), .C(n624), .Y(n4969) );
  NAND2X1 U1138 ( .A(ram[532]), .B(n13002), .Y(n624) );
  OAI21X1 U1139 ( .A(n12744), .B(n13002), .C(n625), .Y(n4970) );
  NAND2X1 U1140 ( .A(ram[533]), .B(n13002), .Y(n625) );
  OAI21X1 U1141 ( .A(n12738), .B(n13002), .C(n626), .Y(n4971) );
  NAND2X1 U1142 ( .A(ram[534]), .B(n13002), .Y(n626) );
  OAI21X1 U1143 ( .A(n12732), .B(n13002), .C(n627), .Y(n4972) );
  NAND2X1 U1144 ( .A(ram[535]), .B(n13002), .Y(n627) );
  OAI21X1 U1145 ( .A(n12726), .B(n13002), .C(n628), .Y(n4973) );
  NAND2X1 U1146 ( .A(ram[536]), .B(n13002), .Y(n628) );
  OAI21X1 U1147 ( .A(n12720), .B(n13002), .C(n629), .Y(n4974) );
  NAND2X1 U1148 ( .A(ram[537]), .B(n13002), .Y(n629) );
  OAI21X1 U1149 ( .A(n12714), .B(n13002), .C(n630), .Y(n4975) );
  NAND2X1 U1150 ( .A(ram[538]), .B(n13002), .Y(n630) );
  OAI21X1 U1151 ( .A(n12708), .B(n13002), .C(n631), .Y(n4976) );
  NAND2X1 U1152 ( .A(ram[539]), .B(n13002), .Y(n631) );
  OAI21X1 U1153 ( .A(n12702), .B(n13002), .C(n632), .Y(n4977) );
  NAND2X1 U1154 ( .A(ram[540]), .B(n13002), .Y(n632) );
  OAI21X1 U1155 ( .A(n12696), .B(n13002), .C(n633), .Y(n4978) );
  NAND2X1 U1156 ( .A(ram[541]), .B(n13002), .Y(n633) );
  OAI21X1 U1157 ( .A(n12690), .B(n13002), .C(n634), .Y(n4979) );
  NAND2X1 U1158 ( .A(ram[542]), .B(n13002), .Y(n634) );
  OAI21X1 U1159 ( .A(n12684), .B(n13002), .C(n635), .Y(n4980) );
  NAND2X1 U1160 ( .A(ram[543]), .B(n13002), .Y(n635) );
  OAI21X1 U1162 ( .A(n12775), .B(n13001), .C(n637), .Y(n4981) );
  NAND2X1 U1163 ( .A(ram[544]), .B(n13001), .Y(n637) );
  OAI21X1 U1164 ( .A(n12769), .B(n13001), .C(n638), .Y(n4982) );
  NAND2X1 U1165 ( .A(ram[545]), .B(n13001), .Y(n638) );
  OAI21X1 U1166 ( .A(n12762), .B(n13001), .C(n639), .Y(n4983) );
  NAND2X1 U1167 ( .A(ram[546]), .B(n13001), .Y(n639) );
  OAI21X1 U1168 ( .A(n12756), .B(n13001), .C(n640), .Y(n4984) );
  NAND2X1 U1169 ( .A(ram[547]), .B(n13001), .Y(n640) );
  OAI21X1 U1170 ( .A(n12750), .B(n13001), .C(n641), .Y(n4985) );
  NAND2X1 U1171 ( .A(ram[548]), .B(n13001), .Y(n641) );
  OAI21X1 U1172 ( .A(n12744), .B(n13001), .C(n642), .Y(n4986) );
  NAND2X1 U1173 ( .A(ram[549]), .B(n13001), .Y(n642) );
  OAI21X1 U1174 ( .A(n12738), .B(n13001), .C(n643), .Y(n4987) );
  NAND2X1 U1175 ( .A(ram[550]), .B(n13001), .Y(n643) );
  OAI21X1 U1176 ( .A(n12732), .B(n13001), .C(n644), .Y(n4988) );
  NAND2X1 U1177 ( .A(ram[551]), .B(n13001), .Y(n644) );
  OAI21X1 U1178 ( .A(n12726), .B(n13001), .C(n645), .Y(n4989) );
  NAND2X1 U1179 ( .A(ram[552]), .B(n13001), .Y(n645) );
  OAI21X1 U1180 ( .A(n12720), .B(n13001), .C(n646), .Y(n4990) );
  NAND2X1 U1181 ( .A(ram[553]), .B(n13001), .Y(n646) );
  OAI21X1 U1182 ( .A(n12714), .B(n13001), .C(n647), .Y(n4991) );
  NAND2X1 U1183 ( .A(ram[554]), .B(n13001), .Y(n647) );
  OAI21X1 U1184 ( .A(n12708), .B(n13001), .C(n648), .Y(n4992) );
  NAND2X1 U1185 ( .A(ram[555]), .B(n13001), .Y(n648) );
  OAI21X1 U1186 ( .A(n12702), .B(n13001), .C(n649), .Y(n4993) );
  NAND2X1 U1187 ( .A(ram[556]), .B(n13001), .Y(n649) );
  OAI21X1 U1188 ( .A(n12696), .B(n13001), .C(n650), .Y(n4994) );
  NAND2X1 U1189 ( .A(ram[557]), .B(n13001), .Y(n650) );
  OAI21X1 U1190 ( .A(n12691), .B(n13001), .C(n651), .Y(n4995) );
  NAND2X1 U1191 ( .A(ram[558]), .B(n13001), .Y(n651) );
  OAI21X1 U1192 ( .A(n12685), .B(n13001), .C(n652), .Y(n4996) );
  NAND2X1 U1193 ( .A(ram[559]), .B(n13001), .Y(n652) );
  OAI21X1 U1195 ( .A(n12774), .B(n13000), .C(n654), .Y(n4997) );
  NAND2X1 U1196 ( .A(ram[560]), .B(n13000), .Y(n654) );
  OAI21X1 U1197 ( .A(n12768), .B(n13000), .C(n655), .Y(n4998) );
  NAND2X1 U1198 ( .A(ram[561]), .B(n13000), .Y(n655) );
  OAI21X1 U1199 ( .A(n12763), .B(n13000), .C(n656), .Y(n4999) );
  NAND2X1 U1200 ( .A(ram[562]), .B(n13000), .Y(n656) );
  OAI21X1 U1201 ( .A(n12757), .B(n13000), .C(n657), .Y(n5000) );
  NAND2X1 U1202 ( .A(ram[563]), .B(n13000), .Y(n657) );
  OAI21X1 U1203 ( .A(n12751), .B(n13000), .C(n658), .Y(n5001) );
  NAND2X1 U1204 ( .A(ram[564]), .B(n13000), .Y(n658) );
  OAI21X1 U1205 ( .A(n12745), .B(n13000), .C(n659), .Y(n5002) );
  NAND2X1 U1206 ( .A(ram[565]), .B(n13000), .Y(n659) );
  OAI21X1 U1207 ( .A(n12739), .B(n13000), .C(n660), .Y(n5003) );
  NAND2X1 U1208 ( .A(ram[566]), .B(n13000), .Y(n660) );
  OAI21X1 U1209 ( .A(n12733), .B(n13000), .C(n661), .Y(n5004) );
  NAND2X1 U1210 ( .A(ram[567]), .B(n13000), .Y(n661) );
  OAI21X1 U1211 ( .A(n12727), .B(n13000), .C(n662), .Y(n5005) );
  NAND2X1 U1212 ( .A(ram[568]), .B(n13000), .Y(n662) );
  OAI21X1 U1213 ( .A(n12721), .B(n13000), .C(n663), .Y(n5006) );
  NAND2X1 U1214 ( .A(ram[569]), .B(n13000), .Y(n663) );
  OAI21X1 U1215 ( .A(n12715), .B(n13000), .C(n664), .Y(n5007) );
  NAND2X1 U1216 ( .A(ram[570]), .B(n13000), .Y(n664) );
  OAI21X1 U1217 ( .A(n12709), .B(n13000), .C(n665), .Y(n5008) );
  NAND2X1 U1218 ( .A(ram[571]), .B(n13000), .Y(n665) );
  OAI21X1 U1219 ( .A(n12703), .B(n13000), .C(n666), .Y(n5009) );
  NAND2X1 U1220 ( .A(ram[572]), .B(n13000), .Y(n666) );
  OAI21X1 U1221 ( .A(n12697), .B(n13000), .C(n667), .Y(n5010) );
  NAND2X1 U1222 ( .A(ram[573]), .B(n13000), .Y(n667) );
  OAI21X1 U1223 ( .A(n12690), .B(n13000), .C(n668), .Y(n5011) );
  NAND2X1 U1224 ( .A(ram[574]), .B(n13000), .Y(n668) );
  OAI21X1 U1225 ( .A(n12684), .B(n13000), .C(n669), .Y(n5012) );
  NAND2X1 U1226 ( .A(ram[575]), .B(n13000), .Y(n669) );
  OAI21X1 U1228 ( .A(n12775), .B(n12999), .C(n671), .Y(n5013) );
  NAND2X1 U1229 ( .A(ram[576]), .B(n12999), .Y(n671) );
  OAI21X1 U1230 ( .A(n12769), .B(n12999), .C(n672), .Y(n5014) );
  NAND2X1 U1231 ( .A(ram[577]), .B(n12999), .Y(n672) );
  OAI21X1 U1232 ( .A(n12762), .B(n12999), .C(n673), .Y(n5015) );
  NAND2X1 U1233 ( .A(ram[578]), .B(n12999), .Y(n673) );
  OAI21X1 U1234 ( .A(n12756), .B(n12999), .C(n674), .Y(n5016) );
  NAND2X1 U1235 ( .A(ram[579]), .B(n12999), .Y(n674) );
  OAI21X1 U1236 ( .A(n12750), .B(n12999), .C(n675), .Y(n5017) );
  NAND2X1 U1237 ( .A(ram[580]), .B(n12999), .Y(n675) );
  OAI21X1 U1238 ( .A(n12744), .B(n12999), .C(n676), .Y(n5018) );
  NAND2X1 U1239 ( .A(ram[581]), .B(n12999), .Y(n676) );
  OAI21X1 U1240 ( .A(n12738), .B(n12999), .C(n677), .Y(n5019) );
  NAND2X1 U1241 ( .A(ram[582]), .B(n12999), .Y(n677) );
  OAI21X1 U1242 ( .A(n12732), .B(n12999), .C(n678), .Y(n5020) );
  NAND2X1 U1243 ( .A(ram[583]), .B(n12999), .Y(n678) );
  OAI21X1 U1244 ( .A(n12726), .B(n12999), .C(n679), .Y(n5021) );
  NAND2X1 U1245 ( .A(ram[584]), .B(n12999), .Y(n679) );
  OAI21X1 U1246 ( .A(n12720), .B(n12999), .C(n680), .Y(n5022) );
  NAND2X1 U1247 ( .A(ram[585]), .B(n12999), .Y(n680) );
  OAI21X1 U1248 ( .A(n12714), .B(n12999), .C(n681), .Y(n5023) );
  NAND2X1 U1249 ( .A(ram[586]), .B(n12999), .Y(n681) );
  OAI21X1 U1250 ( .A(n12708), .B(n12999), .C(n682), .Y(n5024) );
  NAND2X1 U1251 ( .A(ram[587]), .B(n12999), .Y(n682) );
  OAI21X1 U1252 ( .A(n12702), .B(n12999), .C(n683), .Y(n5025) );
  NAND2X1 U1253 ( .A(ram[588]), .B(n12999), .Y(n683) );
  OAI21X1 U1254 ( .A(n12696), .B(n12999), .C(n684), .Y(n5026) );
  NAND2X1 U1255 ( .A(ram[589]), .B(n12999), .Y(n684) );
  OAI21X1 U1256 ( .A(n12691), .B(n12999), .C(n685), .Y(n5027) );
  NAND2X1 U1257 ( .A(ram[590]), .B(n12999), .Y(n685) );
  OAI21X1 U1258 ( .A(n12685), .B(n12999), .C(n686), .Y(n5028) );
  NAND2X1 U1259 ( .A(ram[591]), .B(n12999), .Y(n686) );
  OAI21X1 U1261 ( .A(n12776), .B(n12998), .C(n688), .Y(n5029) );
  NAND2X1 U1262 ( .A(ram[592]), .B(n12998), .Y(n688) );
  OAI21X1 U1263 ( .A(n12770), .B(n12998), .C(n689), .Y(n5030) );
  NAND2X1 U1264 ( .A(ram[593]), .B(n12998), .Y(n689) );
  OAI21X1 U1265 ( .A(n12763), .B(n12998), .C(n690), .Y(n5031) );
  NAND2X1 U1266 ( .A(ram[594]), .B(n12998), .Y(n690) );
  OAI21X1 U1267 ( .A(n12757), .B(n12998), .C(n691), .Y(n5032) );
  NAND2X1 U1268 ( .A(ram[595]), .B(n12998), .Y(n691) );
  OAI21X1 U1269 ( .A(n12751), .B(n12998), .C(n692), .Y(n5033) );
  NAND2X1 U1270 ( .A(ram[596]), .B(n12998), .Y(n692) );
  OAI21X1 U1271 ( .A(n12745), .B(n12998), .C(n693), .Y(n5034) );
  NAND2X1 U1272 ( .A(ram[597]), .B(n12998), .Y(n693) );
  OAI21X1 U1273 ( .A(n12739), .B(n12998), .C(n694), .Y(n5035) );
  NAND2X1 U1274 ( .A(ram[598]), .B(n12998), .Y(n694) );
  OAI21X1 U1275 ( .A(n12733), .B(n12998), .C(n695), .Y(n5036) );
  NAND2X1 U1276 ( .A(ram[599]), .B(n12998), .Y(n695) );
  OAI21X1 U1277 ( .A(n12727), .B(n12998), .C(n696), .Y(n5037) );
  NAND2X1 U1278 ( .A(ram[600]), .B(n12998), .Y(n696) );
  OAI21X1 U1279 ( .A(n12721), .B(n12998), .C(n697), .Y(n5038) );
  NAND2X1 U1280 ( .A(ram[601]), .B(n12998), .Y(n697) );
  OAI21X1 U1281 ( .A(n12715), .B(n12998), .C(n698), .Y(n5039) );
  NAND2X1 U1282 ( .A(ram[602]), .B(n12998), .Y(n698) );
  OAI21X1 U1283 ( .A(n12709), .B(n12998), .C(n699), .Y(n5040) );
  NAND2X1 U1284 ( .A(ram[603]), .B(n12998), .Y(n699) );
  OAI21X1 U1285 ( .A(n12703), .B(n12998), .C(n700), .Y(n5041) );
  NAND2X1 U1286 ( .A(ram[604]), .B(n12998), .Y(n700) );
  OAI21X1 U1287 ( .A(n12697), .B(n12998), .C(n701), .Y(n5042) );
  NAND2X1 U1288 ( .A(ram[605]), .B(n12998), .Y(n701) );
  OAI21X1 U1289 ( .A(n12692), .B(n12998), .C(n702), .Y(n5043) );
  NAND2X1 U1290 ( .A(ram[606]), .B(n12998), .Y(n702) );
  OAI21X1 U1291 ( .A(n12686), .B(n12998), .C(n703), .Y(n5044) );
  NAND2X1 U1292 ( .A(ram[607]), .B(n12998), .Y(n703) );
  OAI21X1 U1294 ( .A(n12775), .B(n12997), .C(n705), .Y(n5045) );
  NAND2X1 U1295 ( .A(ram[608]), .B(n12997), .Y(n705) );
  OAI21X1 U1296 ( .A(n12769), .B(n12997), .C(n706), .Y(n5046) );
  NAND2X1 U1297 ( .A(ram[609]), .B(n12997), .Y(n706) );
  OAI21X1 U1298 ( .A(n12767), .B(n12997), .C(n707), .Y(n5047) );
  NAND2X1 U1299 ( .A(ram[610]), .B(n12997), .Y(n707) );
  OAI21X1 U1300 ( .A(n12761), .B(n12997), .C(n708), .Y(n5048) );
  NAND2X1 U1301 ( .A(ram[611]), .B(n12997), .Y(n708) );
  OAI21X1 U1302 ( .A(n12755), .B(n12997), .C(n709), .Y(n5049) );
  NAND2X1 U1303 ( .A(ram[612]), .B(n12997), .Y(n709) );
  OAI21X1 U1304 ( .A(n12749), .B(n12997), .C(n710), .Y(n5050) );
  NAND2X1 U1305 ( .A(ram[613]), .B(n12997), .Y(n710) );
  OAI21X1 U1306 ( .A(n12743), .B(n12997), .C(n711), .Y(n5051) );
  NAND2X1 U1307 ( .A(ram[614]), .B(n12997), .Y(n711) );
  OAI21X1 U1308 ( .A(n12737), .B(n12997), .C(n712), .Y(n5052) );
  NAND2X1 U1309 ( .A(ram[615]), .B(n12997), .Y(n712) );
  OAI21X1 U1310 ( .A(n12731), .B(n12997), .C(n713), .Y(n5053) );
  NAND2X1 U1311 ( .A(ram[616]), .B(n12997), .Y(n713) );
  OAI21X1 U1312 ( .A(n12725), .B(n12997), .C(n714), .Y(n5054) );
  NAND2X1 U1313 ( .A(ram[617]), .B(n12997), .Y(n714) );
  OAI21X1 U1314 ( .A(n12719), .B(n12997), .C(n715), .Y(n5055) );
  NAND2X1 U1315 ( .A(ram[618]), .B(n12997), .Y(n715) );
  OAI21X1 U1316 ( .A(n12713), .B(n12997), .C(n716), .Y(n5056) );
  NAND2X1 U1317 ( .A(ram[619]), .B(n12997), .Y(n716) );
  OAI21X1 U1318 ( .A(n12707), .B(n12997), .C(n717), .Y(n5057) );
  NAND2X1 U1319 ( .A(ram[620]), .B(n12997), .Y(n717) );
  OAI21X1 U1320 ( .A(n12701), .B(n12997), .C(n718), .Y(n5058) );
  NAND2X1 U1321 ( .A(ram[621]), .B(n12997), .Y(n718) );
  OAI21X1 U1322 ( .A(n12691), .B(n12997), .C(n719), .Y(n5059) );
  NAND2X1 U1323 ( .A(ram[622]), .B(n12997), .Y(n719) );
  OAI21X1 U1324 ( .A(n12685), .B(n12997), .C(n720), .Y(n5060) );
  NAND2X1 U1325 ( .A(ram[623]), .B(n12997), .Y(n720) );
  OAI21X1 U1327 ( .A(n13071), .B(n12996), .C(n722), .Y(n5061) );
  NAND2X1 U1328 ( .A(ram[624]), .B(n12996), .Y(n722) );
  OAI21X1 U1329 ( .A(n13070), .B(n12996), .C(n723), .Y(n5062) );
  NAND2X1 U1330 ( .A(ram[625]), .B(n12996), .Y(n723) );
  OAI21X1 U1331 ( .A(n13069), .B(n12996), .C(n724), .Y(n5063) );
  NAND2X1 U1332 ( .A(ram[626]), .B(n12996), .Y(n724) );
  OAI21X1 U1333 ( .A(n13068), .B(n12996), .C(n725), .Y(n5064) );
  NAND2X1 U1334 ( .A(ram[627]), .B(n12996), .Y(n725) );
  OAI21X1 U1335 ( .A(n13067), .B(n12996), .C(n726), .Y(n5065) );
  NAND2X1 U1336 ( .A(ram[628]), .B(n12996), .Y(n726) );
  OAI21X1 U1337 ( .A(n13066), .B(n12996), .C(n727), .Y(n5066) );
  NAND2X1 U1338 ( .A(ram[629]), .B(n12996), .Y(n727) );
  OAI21X1 U1339 ( .A(n13065), .B(n12996), .C(n728), .Y(n5067) );
  NAND2X1 U1340 ( .A(ram[630]), .B(n12996), .Y(n728) );
  OAI21X1 U1341 ( .A(n13064), .B(n12996), .C(n729), .Y(n5068) );
  NAND2X1 U1342 ( .A(ram[631]), .B(n12996), .Y(n729) );
  OAI21X1 U1343 ( .A(n13063), .B(n12996), .C(n730), .Y(n5069) );
  NAND2X1 U1344 ( .A(ram[632]), .B(n12996), .Y(n730) );
  OAI21X1 U1345 ( .A(n13062), .B(n12996), .C(n731), .Y(n5070) );
  NAND2X1 U1346 ( .A(ram[633]), .B(n12996), .Y(n731) );
  OAI21X1 U1347 ( .A(n13061), .B(n12996), .C(n732), .Y(n5071) );
  NAND2X1 U1348 ( .A(ram[634]), .B(n12996), .Y(n732) );
  OAI21X1 U1349 ( .A(n13060), .B(n12996), .C(n733), .Y(n5072) );
  NAND2X1 U1350 ( .A(ram[635]), .B(n12996), .Y(n733) );
  OAI21X1 U1351 ( .A(n13059), .B(n12996), .C(n734), .Y(n5073) );
  NAND2X1 U1352 ( .A(ram[636]), .B(n12996), .Y(n734) );
  OAI21X1 U1353 ( .A(n13058), .B(n12996), .C(n735), .Y(n5074) );
  NAND2X1 U1354 ( .A(ram[637]), .B(n12996), .Y(n735) );
  OAI21X1 U1355 ( .A(n13057), .B(n12996), .C(n736), .Y(n5075) );
  NAND2X1 U1356 ( .A(ram[638]), .B(n12996), .Y(n736) );
  OAI21X1 U1357 ( .A(n13056), .B(n12996), .C(n737), .Y(n5076) );
  NAND2X1 U1358 ( .A(ram[639]), .B(n12996), .Y(n737) );
  OAI21X1 U1360 ( .A(n13071), .B(n12995), .C(n739), .Y(n5077) );
  NAND2X1 U1361 ( .A(ram[640]), .B(n12995), .Y(n739) );
  OAI21X1 U1362 ( .A(n13070), .B(n12995), .C(n740), .Y(n5078) );
  NAND2X1 U1363 ( .A(ram[641]), .B(n12995), .Y(n740) );
  OAI21X1 U1364 ( .A(n13069), .B(n12995), .C(n741), .Y(n5079) );
  NAND2X1 U1365 ( .A(ram[642]), .B(n12995), .Y(n741) );
  OAI21X1 U1366 ( .A(n13068), .B(n12995), .C(n742), .Y(n5080) );
  NAND2X1 U1367 ( .A(ram[643]), .B(n12995), .Y(n742) );
  OAI21X1 U1368 ( .A(n13067), .B(n12995), .C(n743), .Y(n5081) );
  NAND2X1 U1369 ( .A(ram[644]), .B(n12995), .Y(n743) );
  OAI21X1 U1370 ( .A(n13066), .B(n12995), .C(n744), .Y(n5082) );
  NAND2X1 U1371 ( .A(ram[645]), .B(n12995), .Y(n744) );
  OAI21X1 U1372 ( .A(n13065), .B(n12995), .C(n745), .Y(n5083) );
  NAND2X1 U1373 ( .A(ram[646]), .B(n12995), .Y(n745) );
  OAI21X1 U1374 ( .A(n13064), .B(n12995), .C(n746), .Y(n5084) );
  NAND2X1 U1375 ( .A(ram[647]), .B(n12995), .Y(n746) );
  OAI21X1 U1376 ( .A(n13063), .B(n12995), .C(n747), .Y(n5085) );
  NAND2X1 U1377 ( .A(ram[648]), .B(n12995), .Y(n747) );
  OAI21X1 U1378 ( .A(n13062), .B(n12995), .C(n748), .Y(n5086) );
  NAND2X1 U1379 ( .A(ram[649]), .B(n12995), .Y(n748) );
  OAI21X1 U1380 ( .A(n13061), .B(n12995), .C(n749), .Y(n5087) );
  NAND2X1 U1381 ( .A(ram[650]), .B(n12995), .Y(n749) );
  OAI21X1 U1382 ( .A(n13060), .B(n12995), .C(n750), .Y(n5088) );
  NAND2X1 U1383 ( .A(ram[651]), .B(n12995), .Y(n750) );
  OAI21X1 U1384 ( .A(n13059), .B(n12995), .C(n751), .Y(n5089) );
  NAND2X1 U1385 ( .A(ram[652]), .B(n12995), .Y(n751) );
  OAI21X1 U1386 ( .A(n13058), .B(n12995), .C(n752), .Y(n5090) );
  NAND2X1 U1387 ( .A(ram[653]), .B(n12995), .Y(n752) );
  OAI21X1 U1388 ( .A(n13057), .B(n12995), .C(n753), .Y(n5091) );
  NAND2X1 U1389 ( .A(ram[654]), .B(n12995), .Y(n753) );
  OAI21X1 U1390 ( .A(n13056), .B(n12995), .C(n754), .Y(n5092) );
  NAND2X1 U1391 ( .A(ram[655]), .B(n12995), .Y(n754) );
  OAI21X1 U1393 ( .A(n13071), .B(n12994), .C(n756), .Y(n5093) );
  NAND2X1 U1394 ( .A(ram[656]), .B(n12994), .Y(n756) );
  OAI21X1 U1395 ( .A(n13070), .B(n12994), .C(n757), .Y(n5094) );
  NAND2X1 U1396 ( .A(ram[657]), .B(n12994), .Y(n757) );
  OAI21X1 U1397 ( .A(n13069), .B(n12994), .C(n758), .Y(n5095) );
  NAND2X1 U1398 ( .A(ram[658]), .B(n12994), .Y(n758) );
  OAI21X1 U1399 ( .A(n13068), .B(n12994), .C(n759), .Y(n5096) );
  NAND2X1 U1400 ( .A(ram[659]), .B(n12994), .Y(n759) );
  OAI21X1 U1401 ( .A(n13067), .B(n12994), .C(n760), .Y(n5097) );
  NAND2X1 U1402 ( .A(ram[660]), .B(n12994), .Y(n760) );
  OAI21X1 U1403 ( .A(n13066), .B(n12994), .C(n761), .Y(n5098) );
  NAND2X1 U1404 ( .A(ram[661]), .B(n12994), .Y(n761) );
  OAI21X1 U1405 ( .A(n13065), .B(n12994), .C(n762), .Y(n5099) );
  NAND2X1 U1406 ( .A(ram[662]), .B(n12994), .Y(n762) );
  OAI21X1 U1407 ( .A(n13064), .B(n12994), .C(n763), .Y(n5100) );
  NAND2X1 U1408 ( .A(ram[663]), .B(n12994), .Y(n763) );
  OAI21X1 U1409 ( .A(n13063), .B(n12994), .C(n764), .Y(n5101) );
  NAND2X1 U1410 ( .A(ram[664]), .B(n12994), .Y(n764) );
  OAI21X1 U1411 ( .A(n13062), .B(n12994), .C(n765), .Y(n5102) );
  NAND2X1 U1412 ( .A(ram[665]), .B(n12994), .Y(n765) );
  OAI21X1 U1413 ( .A(n13061), .B(n12994), .C(n766), .Y(n5103) );
  NAND2X1 U1414 ( .A(ram[666]), .B(n12994), .Y(n766) );
  OAI21X1 U1415 ( .A(n13060), .B(n12994), .C(n767), .Y(n5104) );
  NAND2X1 U1416 ( .A(ram[667]), .B(n12994), .Y(n767) );
  OAI21X1 U1417 ( .A(n13059), .B(n12994), .C(n768), .Y(n5105) );
  NAND2X1 U1418 ( .A(ram[668]), .B(n12994), .Y(n768) );
  OAI21X1 U1419 ( .A(n13058), .B(n12994), .C(n769), .Y(n5106) );
  NAND2X1 U1420 ( .A(ram[669]), .B(n12994), .Y(n769) );
  OAI21X1 U1421 ( .A(n13057), .B(n12994), .C(n770), .Y(n5107) );
  NAND2X1 U1422 ( .A(ram[670]), .B(n12994), .Y(n770) );
  OAI21X1 U1423 ( .A(n13056), .B(n12994), .C(n771), .Y(n5108) );
  NAND2X1 U1424 ( .A(ram[671]), .B(n12994), .Y(n771) );
  OAI21X1 U1426 ( .A(n13071), .B(n12993), .C(n773), .Y(n5109) );
  NAND2X1 U1427 ( .A(ram[672]), .B(n12993), .Y(n773) );
  OAI21X1 U1428 ( .A(n13070), .B(n12993), .C(n774), .Y(n5110) );
  NAND2X1 U1429 ( .A(ram[673]), .B(n12993), .Y(n774) );
  OAI21X1 U1430 ( .A(n13069), .B(n12993), .C(n775), .Y(n5111) );
  NAND2X1 U1431 ( .A(ram[674]), .B(n12993), .Y(n775) );
  OAI21X1 U1432 ( .A(n13068), .B(n12993), .C(n776), .Y(n5112) );
  NAND2X1 U1433 ( .A(ram[675]), .B(n12993), .Y(n776) );
  OAI21X1 U1434 ( .A(n13067), .B(n12993), .C(n777), .Y(n5113) );
  NAND2X1 U1435 ( .A(ram[676]), .B(n12993), .Y(n777) );
  OAI21X1 U1436 ( .A(n13066), .B(n12993), .C(n778), .Y(n5114) );
  NAND2X1 U1437 ( .A(ram[677]), .B(n12993), .Y(n778) );
  OAI21X1 U1438 ( .A(n13065), .B(n12993), .C(n779), .Y(n5115) );
  NAND2X1 U1439 ( .A(ram[678]), .B(n12993), .Y(n779) );
  OAI21X1 U1440 ( .A(n13064), .B(n12993), .C(n780), .Y(n5116) );
  NAND2X1 U1441 ( .A(ram[679]), .B(n12993), .Y(n780) );
  OAI21X1 U1442 ( .A(n13063), .B(n12993), .C(n781), .Y(n5117) );
  NAND2X1 U1443 ( .A(ram[680]), .B(n12993), .Y(n781) );
  OAI21X1 U1444 ( .A(n13062), .B(n12993), .C(n782), .Y(n5118) );
  NAND2X1 U1445 ( .A(ram[681]), .B(n12993), .Y(n782) );
  OAI21X1 U1446 ( .A(n13061), .B(n12993), .C(n783), .Y(n5119) );
  NAND2X1 U1447 ( .A(ram[682]), .B(n12993), .Y(n783) );
  OAI21X1 U1448 ( .A(n13060), .B(n12993), .C(n784), .Y(n5120) );
  NAND2X1 U1449 ( .A(ram[683]), .B(n12993), .Y(n784) );
  OAI21X1 U1450 ( .A(n13059), .B(n12993), .C(n785), .Y(n5121) );
  NAND2X1 U1451 ( .A(ram[684]), .B(n12993), .Y(n785) );
  OAI21X1 U1452 ( .A(n13058), .B(n12993), .C(n786), .Y(n5122) );
  NAND2X1 U1453 ( .A(ram[685]), .B(n12993), .Y(n786) );
  OAI21X1 U1454 ( .A(n13057), .B(n12993), .C(n787), .Y(n5123) );
  NAND2X1 U1455 ( .A(ram[686]), .B(n12993), .Y(n787) );
  OAI21X1 U1456 ( .A(n13056), .B(n12993), .C(n788), .Y(n5124) );
  NAND2X1 U1457 ( .A(ram[687]), .B(n12993), .Y(n788) );
  OAI21X1 U1459 ( .A(n13071), .B(n12992), .C(n790), .Y(n5125) );
  NAND2X1 U1460 ( .A(ram[688]), .B(n12992), .Y(n790) );
  OAI21X1 U1461 ( .A(n13070), .B(n12992), .C(n791), .Y(n5126) );
  NAND2X1 U1462 ( .A(ram[689]), .B(n12992), .Y(n791) );
  OAI21X1 U1463 ( .A(n13069), .B(n12992), .C(n792), .Y(n5127) );
  NAND2X1 U1464 ( .A(ram[690]), .B(n12992), .Y(n792) );
  OAI21X1 U1465 ( .A(n13068), .B(n12992), .C(n793), .Y(n5128) );
  NAND2X1 U1466 ( .A(ram[691]), .B(n12992), .Y(n793) );
  OAI21X1 U1467 ( .A(n13067), .B(n12992), .C(n794), .Y(n5129) );
  NAND2X1 U1468 ( .A(ram[692]), .B(n12992), .Y(n794) );
  OAI21X1 U1469 ( .A(n13066), .B(n12992), .C(n795), .Y(n5130) );
  NAND2X1 U1470 ( .A(ram[693]), .B(n12992), .Y(n795) );
  OAI21X1 U1471 ( .A(n13065), .B(n12992), .C(n796), .Y(n5131) );
  NAND2X1 U1472 ( .A(ram[694]), .B(n12992), .Y(n796) );
  OAI21X1 U1473 ( .A(n13064), .B(n12992), .C(n797), .Y(n5132) );
  NAND2X1 U1474 ( .A(ram[695]), .B(n12992), .Y(n797) );
  OAI21X1 U1475 ( .A(n13063), .B(n12992), .C(n798), .Y(n5133) );
  NAND2X1 U1476 ( .A(ram[696]), .B(n12992), .Y(n798) );
  OAI21X1 U1477 ( .A(n13062), .B(n12992), .C(n799), .Y(n5134) );
  NAND2X1 U1478 ( .A(ram[697]), .B(n12992), .Y(n799) );
  OAI21X1 U1479 ( .A(n13061), .B(n12992), .C(n800), .Y(n5135) );
  NAND2X1 U1480 ( .A(ram[698]), .B(n12992), .Y(n800) );
  OAI21X1 U1481 ( .A(n13060), .B(n12992), .C(n801), .Y(n5136) );
  NAND2X1 U1482 ( .A(ram[699]), .B(n12992), .Y(n801) );
  OAI21X1 U1483 ( .A(n13059), .B(n12992), .C(n802), .Y(n5137) );
  NAND2X1 U1484 ( .A(ram[700]), .B(n12992), .Y(n802) );
  OAI21X1 U1485 ( .A(n13058), .B(n12992), .C(n803), .Y(n5138) );
  NAND2X1 U1486 ( .A(ram[701]), .B(n12992), .Y(n803) );
  OAI21X1 U1487 ( .A(n13057), .B(n12992), .C(n804), .Y(n5139) );
  NAND2X1 U1488 ( .A(ram[702]), .B(n12992), .Y(n804) );
  OAI21X1 U1489 ( .A(n13056), .B(n12992), .C(n805), .Y(n5140) );
  NAND2X1 U1490 ( .A(ram[703]), .B(n12992), .Y(n805) );
  OAI21X1 U1492 ( .A(n13071), .B(n12991), .C(n807), .Y(n5141) );
  NAND2X1 U1493 ( .A(ram[704]), .B(n12991), .Y(n807) );
  OAI21X1 U1494 ( .A(n13070), .B(n12991), .C(n808), .Y(n5142) );
  NAND2X1 U1495 ( .A(ram[705]), .B(n12991), .Y(n808) );
  OAI21X1 U1496 ( .A(n13069), .B(n12991), .C(n809), .Y(n5143) );
  NAND2X1 U1497 ( .A(ram[706]), .B(n12991), .Y(n809) );
  OAI21X1 U1498 ( .A(n13068), .B(n12991), .C(n810), .Y(n5144) );
  NAND2X1 U1499 ( .A(ram[707]), .B(n12991), .Y(n810) );
  OAI21X1 U1500 ( .A(n13067), .B(n12991), .C(n811), .Y(n5145) );
  NAND2X1 U1501 ( .A(ram[708]), .B(n12991), .Y(n811) );
  OAI21X1 U1502 ( .A(n13066), .B(n12991), .C(n812), .Y(n5146) );
  NAND2X1 U1503 ( .A(ram[709]), .B(n12991), .Y(n812) );
  OAI21X1 U1504 ( .A(n13065), .B(n12991), .C(n813), .Y(n5147) );
  NAND2X1 U1505 ( .A(ram[710]), .B(n12991), .Y(n813) );
  OAI21X1 U1506 ( .A(n13064), .B(n12991), .C(n814), .Y(n5148) );
  NAND2X1 U1507 ( .A(ram[711]), .B(n12991), .Y(n814) );
  OAI21X1 U1508 ( .A(n13063), .B(n12991), .C(n815), .Y(n5149) );
  NAND2X1 U1509 ( .A(ram[712]), .B(n12991), .Y(n815) );
  OAI21X1 U1510 ( .A(n13062), .B(n12991), .C(n816), .Y(n5150) );
  NAND2X1 U1511 ( .A(ram[713]), .B(n12991), .Y(n816) );
  OAI21X1 U1512 ( .A(n13061), .B(n12991), .C(n817), .Y(n5151) );
  NAND2X1 U1513 ( .A(ram[714]), .B(n12991), .Y(n817) );
  OAI21X1 U1514 ( .A(n13060), .B(n12991), .C(n818), .Y(n5152) );
  NAND2X1 U1515 ( .A(ram[715]), .B(n12991), .Y(n818) );
  OAI21X1 U1516 ( .A(n13059), .B(n12991), .C(n819), .Y(n5153) );
  NAND2X1 U1517 ( .A(ram[716]), .B(n12991), .Y(n819) );
  OAI21X1 U1518 ( .A(n13058), .B(n12991), .C(n820), .Y(n5154) );
  NAND2X1 U1519 ( .A(ram[717]), .B(n12991), .Y(n820) );
  OAI21X1 U1520 ( .A(n13057), .B(n12991), .C(n821), .Y(n5155) );
  NAND2X1 U1521 ( .A(ram[718]), .B(n12991), .Y(n821) );
  OAI21X1 U1522 ( .A(n13056), .B(n12991), .C(n822), .Y(n5156) );
  NAND2X1 U1523 ( .A(ram[719]), .B(n12991), .Y(n822) );
  OAI21X1 U1525 ( .A(n13071), .B(n12990), .C(n824), .Y(n5157) );
  NAND2X1 U1526 ( .A(ram[720]), .B(n12990), .Y(n824) );
  OAI21X1 U1527 ( .A(n13070), .B(n12990), .C(n825), .Y(n5158) );
  NAND2X1 U1528 ( .A(ram[721]), .B(n12990), .Y(n825) );
  OAI21X1 U1529 ( .A(n13069), .B(n12990), .C(n826), .Y(n5159) );
  NAND2X1 U1530 ( .A(ram[722]), .B(n12990), .Y(n826) );
  OAI21X1 U1531 ( .A(n13068), .B(n12990), .C(n827), .Y(n5160) );
  NAND2X1 U1532 ( .A(ram[723]), .B(n12990), .Y(n827) );
  OAI21X1 U1533 ( .A(n13067), .B(n12990), .C(n828), .Y(n5161) );
  NAND2X1 U1534 ( .A(ram[724]), .B(n12990), .Y(n828) );
  OAI21X1 U1535 ( .A(n13066), .B(n12990), .C(n829), .Y(n5162) );
  NAND2X1 U1536 ( .A(ram[725]), .B(n12990), .Y(n829) );
  OAI21X1 U1537 ( .A(n13065), .B(n12990), .C(n830), .Y(n5163) );
  NAND2X1 U1538 ( .A(ram[726]), .B(n12990), .Y(n830) );
  OAI21X1 U1539 ( .A(n13064), .B(n12990), .C(n831), .Y(n5164) );
  NAND2X1 U1540 ( .A(ram[727]), .B(n12990), .Y(n831) );
  OAI21X1 U1541 ( .A(n13063), .B(n12990), .C(n832), .Y(n5165) );
  NAND2X1 U1542 ( .A(ram[728]), .B(n12990), .Y(n832) );
  OAI21X1 U1543 ( .A(n13062), .B(n12990), .C(n833), .Y(n5166) );
  NAND2X1 U1544 ( .A(ram[729]), .B(n12990), .Y(n833) );
  OAI21X1 U1545 ( .A(n13061), .B(n12990), .C(n834), .Y(n5167) );
  NAND2X1 U1546 ( .A(ram[730]), .B(n12990), .Y(n834) );
  OAI21X1 U1547 ( .A(n13060), .B(n12990), .C(n835), .Y(n5168) );
  NAND2X1 U1548 ( .A(ram[731]), .B(n12990), .Y(n835) );
  OAI21X1 U1549 ( .A(n13059), .B(n12990), .C(n836), .Y(n5169) );
  NAND2X1 U1550 ( .A(ram[732]), .B(n12990), .Y(n836) );
  OAI21X1 U1551 ( .A(n13058), .B(n12990), .C(n837), .Y(n5170) );
  NAND2X1 U1552 ( .A(ram[733]), .B(n12990), .Y(n837) );
  OAI21X1 U1553 ( .A(n13057), .B(n12990), .C(n838), .Y(n5171) );
  NAND2X1 U1554 ( .A(ram[734]), .B(n12990), .Y(n838) );
  OAI21X1 U1555 ( .A(n13056), .B(n12990), .C(n839), .Y(n5172) );
  NAND2X1 U1556 ( .A(ram[735]), .B(n12990), .Y(n839) );
  OAI21X1 U1558 ( .A(n13071), .B(n12989), .C(n841), .Y(n5173) );
  NAND2X1 U1559 ( .A(ram[736]), .B(n12989), .Y(n841) );
  OAI21X1 U1560 ( .A(n13070), .B(n12989), .C(n842), .Y(n5174) );
  NAND2X1 U1561 ( .A(ram[737]), .B(n12989), .Y(n842) );
  OAI21X1 U1562 ( .A(n13069), .B(n12989), .C(n843), .Y(n5175) );
  NAND2X1 U1563 ( .A(ram[738]), .B(n12989), .Y(n843) );
  OAI21X1 U1564 ( .A(n13068), .B(n12989), .C(n844), .Y(n5176) );
  NAND2X1 U1565 ( .A(ram[739]), .B(n12989), .Y(n844) );
  OAI21X1 U1566 ( .A(n13067), .B(n12989), .C(n845), .Y(n5177) );
  NAND2X1 U1567 ( .A(ram[740]), .B(n12989), .Y(n845) );
  OAI21X1 U1568 ( .A(n13066), .B(n12989), .C(n846), .Y(n5178) );
  NAND2X1 U1569 ( .A(ram[741]), .B(n12989), .Y(n846) );
  OAI21X1 U1570 ( .A(n13065), .B(n12989), .C(n847), .Y(n5179) );
  NAND2X1 U1571 ( .A(ram[742]), .B(n12989), .Y(n847) );
  OAI21X1 U1572 ( .A(n13064), .B(n12989), .C(n848), .Y(n5180) );
  NAND2X1 U1573 ( .A(ram[743]), .B(n12989), .Y(n848) );
  OAI21X1 U1574 ( .A(n13063), .B(n12989), .C(n849), .Y(n5181) );
  NAND2X1 U1575 ( .A(ram[744]), .B(n12989), .Y(n849) );
  OAI21X1 U1576 ( .A(n13062), .B(n12989), .C(n850), .Y(n5182) );
  NAND2X1 U1577 ( .A(ram[745]), .B(n12989), .Y(n850) );
  OAI21X1 U1578 ( .A(n13061), .B(n12989), .C(n851), .Y(n5183) );
  NAND2X1 U1579 ( .A(ram[746]), .B(n12989), .Y(n851) );
  OAI21X1 U1580 ( .A(n13060), .B(n12989), .C(n852), .Y(n5184) );
  NAND2X1 U1581 ( .A(ram[747]), .B(n12989), .Y(n852) );
  OAI21X1 U1582 ( .A(n13059), .B(n12989), .C(n853), .Y(n5185) );
  NAND2X1 U1583 ( .A(ram[748]), .B(n12989), .Y(n853) );
  OAI21X1 U1584 ( .A(n13058), .B(n12989), .C(n854), .Y(n5186) );
  NAND2X1 U1585 ( .A(ram[749]), .B(n12989), .Y(n854) );
  OAI21X1 U1586 ( .A(n13057), .B(n12989), .C(n855), .Y(n5187) );
  NAND2X1 U1587 ( .A(ram[750]), .B(n12989), .Y(n855) );
  OAI21X1 U1588 ( .A(n13056), .B(n12989), .C(n856), .Y(n5188) );
  NAND2X1 U1589 ( .A(ram[751]), .B(n12989), .Y(n856) );
  OAI21X1 U1591 ( .A(n13071), .B(n12988), .C(n858), .Y(n5189) );
  NAND2X1 U1592 ( .A(ram[752]), .B(n12988), .Y(n858) );
  OAI21X1 U1593 ( .A(n13070), .B(n12988), .C(n859), .Y(n5190) );
  NAND2X1 U1594 ( .A(ram[753]), .B(n12988), .Y(n859) );
  OAI21X1 U1595 ( .A(n13069), .B(n12988), .C(n860), .Y(n5191) );
  NAND2X1 U1596 ( .A(ram[754]), .B(n12988), .Y(n860) );
  OAI21X1 U1597 ( .A(n13068), .B(n12988), .C(n861), .Y(n5192) );
  NAND2X1 U1598 ( .A(ram[755]), .B(n12988), .Y(n861) );
  OAI21X1 U1599 ( .A(n13067), .B(n12988), .C(n862), .Y(n5193) );
  NAND2X1 U1600 ( .A(ram[756]), .B(n12988), .Y(n862) );
  OAI21X1 U1601 ( .A(n13066), .B(n12988), .C(n863), .Y(n5194) );
  NAND2X1 U1602 ( .A(ram[757]), .B(n12988), .Y(n863) );
  OAI21X1 U1603 ( .A(n13065), .B(n12988), .C(n864), .Y(n5195) );
  NAND2X1 U1604 ( .A(ram[758]), .B(n12988), .Y(n864) );
  OAI21X1 U1605 ( .A(n13064), .B(n12988), .C(n865), .Y(n5196) );
  NAND2X1 U1606 ( .A(ram[759]), .B(n12988), .Y(n865) );
  OAI21X1 U1607 ( .A(n13063), .B(n12988), .C(n866), .Y(n5197) );
  NAND2X1 U1608 ( .A(ram[760]), .B(n12988), .Y(n866) );
  OAI21X1 U1609 ( .A(n13062), .B(n12988), .C(n867), .Y(n5198) );
  NAND2X1 U1610 ( .A(ram[761]), .B(n12988), .Y(n867) );
  OAI21X1 U1611 ( .A(n13061), .B(n12988), .C(n868), .Y(n5199) );
  NAND2X1 U1612 ( .A(ram[762]), .B(n12988), .Y(n868) );
  OAI21X1 U1613 ( .A(n13060), .B(n12988), .C(n869), .Y(n5200) );
  NAND2X1 U1614 ( .A(ram[763]), .B(n12988), .Y(n869) );
  OAI21X1 U1615 ( .A(n13059), .B(n12988), .C(n870), .Y(n5201) );
  NAND2X1 U1616 ( .A(ram[764]), .B(n12988), .Y(n870) );
  OAI21X1 U1617 ( .A(n13058), .B(n12988), .C(n871), .Y(n5202) );
  NAND2X1 U1618 ( .A(ram[765]), .B(n12988), .Y(n871) );
  OAI21X1 U1619 ( .A(n13057), .B(n12988), .C(n872), .Y(n5203) );
  NAND2X1 U1620 ( .A(ram[766]), .B(n12988), .Y(n872) );
  OAI21X1 U1621 ( .A(n13056), .B(n12988), .C(n873), .Y(n5204) );
  NAND2X1 U1622 ( .A(ram[767]), .B(n12988), .Y(n873) );
  NAND3X1 U1624 ( .A(mem_write_en), .B(n326), .C(n875), .Y(n874) );
  OAI21X1 U1625 ( .A(n13071), .B(n12987), .C(n877), .Y(n5205) );
  NAND2X1 U1626 ( .A(ram[768]), .B(n12987), .Y(n877) );
  OAI21X1 U1627 ( .A(n13070), .B(n12987), .C(n878), .Y(n5206) );
  NAND2X1 U1628 ( .A(ram[769]), .B(n12987), .Y(n878) );
  OAI21X1 U1629 ( .A(n13069), .B(n12987), .C(n879), .Y(n5207) );
  NAND2X1 U1630 ( .A(ram[770]), .B(n12987), .Y(n879) );
  OAI21X1 U1631 ( .A(n13068), .B(n12987), .C(n880), .Y(n5208) );
  NAND2X1 U1632 ( .A(ram[771]), .B(n12987), .Y(n880) );
  OAI21X1 U1633 ( .A(n13067), .B(n12987), .C(n881), .Y(n5209) );
  NAND2X1 U1634 ( .A(ram[772]), .B(n12987), .Y(n881) );
  OAI21X1 U1635 ( .A(n13066), .B(n12987), .C(n882), .Y(n5210) );
  NAND2X1 U1636 ( .A(ram[773]), .B(n12987), .Y(n882) );
  OAI21X1 U1637 ( .A(n13065), .B(n12987), .C(n883), .Y(n5211) );
  NAND2X1 U1638 ( .A(ram[774]), .B(n12987), .Y(n883) );
  OAI21X1 U1639 ( .A(n13064), .B(n12987), .C(n884), .Y(n5212) );
  NAND2X1 U1640 ( .A(ram[775]), .B(n12987), .Y(n884) );
  OAI21X1 U1641 ( .A(n13063), .B(n12987), .C(n885), .Y(n5213) );
  NAND2X1 U1642 ( .A(ram[776]), .B(n12987), .Y(n885) );
  OAI21X1 U1643 ( .A(n13062), .B(n12987), .C(n886), .Y(n5214) );
  NAND2X1 U1644 ( .A(ram[777]), .B(n12987), .Y(n886) );
  OAI21X1 U1645 ( .A(n13061), .B(n12987), .C(n887), .Y(n5215) );
  NAND2X1 U1646 ( .A(ram[778]), .B(n12987), .Y(n887) );
  OAI21X1 U1647 ( .A(n13060), .B(n12987), .C(n888), .Y(n5216) );
  NAND2X1 U1648 ( .A(ram[779]), .B(n12987), .Y(n888) );
  OAI21X1 U1649 ( .A(n13059), .B(n12987), .C(n889), .Y(n5217) );
  NAND2X1 U1650 ( .A(ram[780]), .B(n12987), .Y(n889) );
  OAI21X1 U1651 ( .A(n13058), .B(n12987), .C(n890), .Y(n5218) );
  NAND2X1 U1652 ( .A(ram[781]), .B(n12987), .Y(n890) );
  OAI21X1 U1653 ( .A(n13057), .B(n12987), .C(n891), .Y(n5219) );
  NAND2X1 U1654 ( .A(ram[782]), .B(n12987), .Y(n891) );
  OAI21X1 U1655 ( .A(n13056), .B(n12987), .C(n892), .Y(n5220) );
  NAND2X1 U1656 ( .A(ram[783]), .B(n12987), .Y(n892) );
  OAI21X1 U1658 ( .A(n13071), .B(n12986), .C(n894), .Y(n5221) );
  NAND2X1 U1659 ( .A(ram[784]), .B(n12986), .Y(n894) );
  OAI21X1 U1660 ( .A(n13070), .B(n12986), .C(n895), .Y(n5222) );
  NAND2X1 U1661 ( .A(ram[785]), .B(n12986), .Y(n895) );
  OAI21X1 U1662 ( .A(n13069), .B(n12986), .C(n896), .Y(n5223) );
  NAND2X1 U1663 ( .A(ram[786]), .B(n12986), .Y(n896) );
  OAI21X1 U1664 ( .A(n13068), .B(n12986), .C(n897), .Y(n5224) );
  NAND2X1 U1665 ( .A(ram[787]), .B(n12986), .Y(n897) );
  OAI21X1 U1666 ( .A(n13067), .B(n12986), .C(n898), .Y(n5225) );
  NAND2X1 U1667 ( .A(ram[788]), .B(n12986), .Y(n898) );
  OAI21X1 U1668 ( .A(n13066), .B(n12986), .C(n899), .Y(n5226) );
  NAND2X1 U1669 ( .A(ram[789]), .B(n12986), .Y(n899) );
  OAI21X1 U1670 ( .A(n13065), .B(n12986), .C(n900), .Y(n5227) );
  NAND2X1 U1671 ( .A(ram[790]), .B(n12986), .Y(n900) );
  OAI21X1 U1672 ( .A(n13064), .B(n12986), .C(n901), .Y(n5228) );
  NAND2X1 U1673 ( .A(ram[791]), .B(n12986), .Y(n901) );
  OAI21X1 U1674 ( .A(n13063), .B(n12986), .C(n902), .Y(n5229) );
  NAND2X1 U1675 ( .A(ram[792]), .B(n12986), .Y(n902) );
  OAI21X1 U1676 ( .A(n13062), .B(n12986), .C(n903), .Y(n5230) );
  NAND2X1 U1677 ( .A(ram[793]), .B(n12986), .Y(n903) );
  OAI21X1 U1678 ( .A(n13061), .B(n12986), .C(n904), .Y(n5231) );
  NAND2X1 U1679 ( .A(ram[794]), .B(n12986), .Y(n904) );
  OAI21X1 U1680 ( .A(n13060), .B(n12986), .C(n905), .Y(n5232) );
  NAND2X1 U1681 ( .A(ram[795]), .B(n12986), .Y(n905) );
  OAI21X1 U1682 ( .A(n13059), .B(n12986), .C(n906), .Y(n5233) );
  NAND2X1 U1683 ( .A(ram[796]), .B(n12986), .Y(n906) );
  OAI21X1 U1684 ( .A(n13058), .B(n12986), .C(n907), .Y(n5234) );
  NAND2X1 U1685 ( .A(ram[797]), .B(n12986), .Y(n907) );
  OAI21X1 U1686 ( .A(n13057), .B(n12986), .C(n908), .Y(n5235) );
  NAND2X1 U1687 ( .A(ram[798]), .B(n12986), .Y(n908) );
  OAI21X1 U1688 ( .A(n13056), .B(n12986), .C(n909), .Y(n5236) );
  NAND2X1 U1689 ( .A(ram[799]), .B(n12986), .Y(n909) );
  OAI21X1 U1691 ( .A(n12774), .B(n12985), .C(n911), .Y(n5237) );
  NAND2X1 U1692 ( .A(ram[800]), .B(n12985), .Y(n911) );
  OAI21X1 U1693 ( .A(n12768), .B(n12985), .C(n912), .Y(n5238) );
  NAND2X1 U1694 ( .A(ram[801]), .B(n12985), .Y(n912) );
  OAI21X1 U1695 ( .A(n13069), .B(n12985), .C(n913), .Y(n5239) );
  NAND2X1 U1696 ( .A(ram[802]), .B(n12985), .Y(n913) );
  OAI21X1 U1697 ( .A(n13068), .B(n12985), .C(n914), .Y(n5240) );
  NAND2X1 U1698 ( .A(ram[803]), .B(n12985), .Y(n914) );
  OAI21X1 U1699 ( .A(n13067), .B(n12985), .C(n915), .Y(n5241) );
  NAND2X1 U1700 ( .A(ram[804]), .B(n12985), .Y(n915) );
  OAI21X1 U1701 ( .A(n13066), .B(n12985), .C(n916), .Y(n5242) );
  NAND2X1 U1702 ( .A(ram[805]), .B(n12985), .Y(n916) );
  OAI21X1 U1703 ( .A(n13065), .B(n12985), .C(n917), .Y(n5243) );
  NAND2X1 U1704 ( .A(ram[806]), .B(n12985), .Y(n917) );
  OAI21X1 U1705 ( .A(n13064), .B(n12985), .C(n918), .Y(n5244) );
  NAND2X1 U1706 ( .A(ram[807]), .B(n12985), .Y(n918) );
  OAI21X1 U1707 ( .A(n13063), .B(n12985), .C(n919), .Y(n5245) );
  NAND2X1 U1708 ( .A(ram[808]), .B(n12985), .Y(n919) );
  OAI21X1 U1709 ( .A(n13062), .B(n12985), .C(n920), .Y(n5246) );
  NAND2X1 U1710 ( .A(ram[809]), .B(n12985), .Y(n920) );
  OAI21X1 U1711 ( .A(n13061), .B(n12985), .C(n921), .Y(n5247) );
  NAND2X1 U1712 ( .A(ram[810]), .B(n12985), .Y(n921) );
  OAI21X1 U1713 ( .A(n13060), .B(n12985), .C(n922), .Y(n5248) );
  NAND2X1 U1714 ( .A(ram[811]), .B(n12985), .Y(n922) );
  OAI21X1 U1715 ( .A(n13059), .B(n12985), .C(n923), .Y(n5249) );
  NAND2X1 U1716 ( .A(ram[812]), .B(n12985), .Y(n923) );
  OAI21X1 U1717 ( .A(n13058), .B(n12985), .C(n924), .Y(n5250) );
  NAND2X1 U1718 ( .A(ram[813]), .B(n12985), .Y(n924) );
  OAI21X1 U1719 ( .A(n12690), .B(n12985), .C(n925), .Y(n5251) );
  NAND2X1 U1720 ( .A(ram[814]), .B(n12985), .Y(n925) );
  OAI21X1 U1721 ( .A(n12684), .B(n12985), .C(n926), .Y(n5252) );
  NAND2X1 U1722 ( .A(ram[815]), .B(n12985), .Y(n926) );
  OAI21X1 U1724 ( .A(n12775), .B(n12984), .C(n928), .Y(n5253) );
  NAND2X1 U1725 ( .A(ram[816]), .B(n12984), .Y(n928) );
  OAI21X1 U1726 ( .A(n12769), .B(n12984), .C(n929), .Y(n5254) );
  NAND2X1 U1727 ( .A(ram[817]), .B(n12984), .Y(n929) );
  OAI21X1 U1728 ( .A(n13069), .B(n12984), .C(n930), .Y(n5255) );
  NAND2X1 U1729 ( .A(ram[818]), .B(n12984), .Y(n930) );
  OAI21X1 U1730 ( .A(n13068), .B(n12984), .C(n931), .Y(n5256) );
  NAND2X1 U1731 ( .A(ram[819]), .B(n12984), .Y(n931) );
  OAI21X1 U1732 ( .A(n13067), .B(n12984), .C(n932), .Y(n5257) );
  NAND2X1 U1733 ( .A(ram[820]), .B(n12984), .Y(n932) );
  OAI21X1 U1734 ( .A(n13066), .B(n12984), .C(n933), .Y(n5258) );
  NAND2X1 U1735 ( .A(ram[821]), .B(n12984), .Y(n933) );
  OAI21X1 U1736 ( .A(n13065), .B(n12984), .C(n934), .Y(n5259) );
  NAND2X1 U1737 ( .A(ram[822]), .B(n12984), .Y(n934) );
  OAI21X1 U1738 ( .A(n13064), .B(n12984), .C(n935), .Y(n5260) );
  NAND2X1 U1739 ( .A(ram[823]), .B(n12984), .Y(n935) );
  OAI21X1 U1740 ( .A(n13063), .B(n12984), .C(n936), .Y(n5261) );
  NAND2X1 U1741 ( .A(ram[824]), .B(n12984), .Y(n936) );
  OAI21X1 U1742 ( .A(n13062), .B(n12984), .C(n937), .Y(n5262) );
  NAND2X1 U1743 ( .A(ram[825]), .B(n12984), .Y(n937) );
  OAI21X1 U1744 ( .A(n13061), .B(n12984), .C(n938), .Y(n5263) );
  NAND2X1 U1745 ( .A(ram[826]), .B(n12984), .Y(n938) );
  OAI21X1 U1746 ( .A(n13060), .B(n12984), .C(n939), .Y(n5264) );
  NAND2X1 U1747 ( .A(ram[827]), .B(n12984), .Y(n939) );
  OAI21X1 U1748 ( .A(n13059), .B(n12984), .C(n940), .Y(n5265) );
  NAND2X1 U1749 ( .A(ram[828]), .B(n12984), .Y(n940) );
  OAI21X1 U1750 ( .A(n13058), .B(n12984), .C(n941), .Y(n5266) );
  NAND2X1 U1751 ( .A(ram[829]), .B(n12984), .Y(n941) );
  OAI21X1 U1752 ( .A(n12691), .B(n12984), .C(n942), .Y(n5267) );
  NAND2X1 U1753 ( .A(ram[830]), .B(n12984), .Y(n942) );
  OAI21X1 U1754 ( .A(n12685), .B(n12984), .C(n943), .Y(n5268) );
  NAND2X1 U1755 ( .A(ram[831]), .B(n12984), .Y(n943) );
  OAI21X1 U1757 ( .A(n13071), .B(n12983), .C(n945), .Y(n5269) );
  NAND2X1 U1758 ( .A(ram[832]), .B(n12983), .Y(n945) );
  OAI21X1 U1759 ( .A(n13070), .B(n12983), .C(n946), .Y(n5270) );
  NAND2X1 U1760 ( .A(ram[833]), .B(n12983), .Y(n946) );
  OAI21X1 U1761 ( .A(n13069), .B(n12983), .C(n947), .Y(n5271) );
  NAND2X1 U1762 ( .A(ram[834]), .B(n12983), .Y(n947) );
  OAI21X1 U1763 ( .A(n13068), .B(n12983), .C(n948), .Y(n5272) );
  NAND2X1 U1764 ( .A(ram[835]), .B(n12983), .Y(n948) );
  OAI21X1 U1765 ( .A(n13067), .B(n12983), .C(n949), .Y(n5273) );
  NAND2X1 U1766 ( .A(ram[836]), .B(n12983), .Y(n949) );
  OAI21X1 U1767 ( .A(n13066), .B(n12983), .C(n950), .Y(n5274) );
  NAND2X1 U1768 ( .A(ram[837]), .B(n12983), .Y(n950) );
  OAI21X1 U1769 ( .A(n13065), .B(n12983), .C(n951), .Y(n5275) );
  NAND2X1 U1770 ( .A(ram[838]), .B(n12983), .Y(n951) );
  OAI21X1 U1771 ( .A(n13064), .B(n12983), .C(n952), .Y(n5276) );
  NAND2X1 U1772 ( .A(ram[839]), .B(n12983), .Y(n952) );
  OAI21X1 U1773 ( .A(n13063), .B(n12983), .C(n953), .Y(n5277) );
  NAND2X1 U1774 ( .A(ram[840]), .B(n12983), .Y(n953) );
  OAI21X1 U1775 ( .A(n13062), .B(n12983), .C(n954), .Y(n5278) );
  NAND2X1 U1776 ( .A(ram[841]), .B(n12983), .Y(n954) );
  OAI21X1 U1777 ( .A(n13061), .B(n12983), .C(n955), .Y(n5279) );
  NAND2X1 U1778 ( .A(ram[842]), .B(n12983), .Y(n955) );
  OAI21X1 U1779 ( .A(n13060), .B(n12983), .C(n956), .Y(n5280) );
  NAND2X1 U1780 ( .A(ram[843]), .B(n12983), .Y(n956) );
  OAI21X1 U1781 ( .A(n13059), .B(n12983), .C(n957), .Y(n5281) );
  NAND2X1 U1782 ( .A(ram[844]), .B(n12983), .Y(n957) );
  OAI21X1 U1783 ( .A(n13058), .B(n12983), .C(n958), .Y(n5282) );
  NAND2X1 U1784 ( .A(ram[845]), .B(n12983), .Y(n958) );
  OAI21X1 U1785 ( .A(n13057), .B(n12983), .C(n959), .Y(n5283) );
  NAND2X1 U1786 ( .A(ram[846]), .B(n12983), .Y(n959) );
  OAI21X1 U1787 ( .A(n13056), .B(n12983), .C(n960), .Y(n5284) );
  NAND2X1 U1788 ( .A(ram[847]), .B(n12983), .Y(n960) );
  OAI21X1 U1790 ( .A(n13071), .B(n12982), .C(n962), .Y(n5285) );
  NAND2X1 U1791 ( .A(ram[848]), .B(n12982), .Y(n962) );
  OAI21X1 U1792 ( .A(n13070), .B(n12982), .C(n963), .Y(n5286) );
  NAND2X1 U1793 ( .A(ram[849]), .B(n12982), .Y(n963) );
  OAI21X1 U1794 ( .A(n13069), .B(n12982), .C(n964), .Y(n5287) );
  NAND2X1 U1795 ( .A(ram[850]), .B(n12982), .Y(n964) );
  OAI21X1 U1796 ( .A(n13068), .B(n12982), .C(n965), .Y(n5288) );
  NAND2X1 U1797 ( .A(ram[851]), .B(n12982), .Y(n965) );
  OAI21X1 U1798 ( .A(n13067), .B(n12982), .C(n966), .Y(n5289) );
  NAND2X1 U1799 ( .A(ram[852]), .B(n12982), .Y(n966) );
  OAI21X1 U1800 ( .A(n13066), .B(n12982), .C(n967), .Y(n5290) );
  NAND2X1 U1801 ( .A(ram[853]), .B(n12982), .Y(n967) );
  OAI21X1 U1802 ( .A(n13065), .B(n12982), .C(n968), .Y(n5291) );
  NAND2X1 U1803 ( .A(ram[854]), .B(n12982), .Y(n968) );
  OAI21X1 U1804 ( .A(n13064), .B(n12982), .C(n969), .Y(n5292) );
  NAND2X1 U1805 ( .A(ram[855]), .B(n12982), .Y(n969) );
  OAI21X1 U1806 ( .A(n13063), .B(n12982), .C(n970), .Y(n5293) );
  NAND2X1 U1807 ( .A(ram[856]), .B(n12982), .Y(n970) );
  OAI21X1 U1808 ( .A(n13062), .B(n12982), .C(n971), .Y(n5294) );
  NAND2X1 U1809 ( .A(ram[857]), .B(n12982), .Y(n971) );
  OAI21X1 U1810 ( .A(n13061), .B(n12982), .C(n972), .Y(n5295) );
  NAND2X1 U1811 ( .A(ram[858]), .B(n12982), .Y(n972) );
  OAI21X1 U1812 ( .A(n13060), .B(n12982), .C(n973), .Y(n5296) );
  NAND2X1 U1813 ( .A(ram[859]), .B(n12982), .Y(n973) );
  OAI21X1 U1814 ( .A(n13059), .B(n12982), .C(n974), .Y(n5297) );
  NAND2X1 U1815 ( .A(ram[860]), .B(n12982), .Y(n974) );
  OAI21X1 U1816 ( .A(n13058), .B(n12982), .C(n975), .Y(n5298) );
  NAND2X1 U1817 ( .A(ram[861]), .B(n12982), .Y(n975) );
  OAI21X1 U1818 ( .A(n13057), .B(n12982), .C(n976), .Y(n5299) );
  NAND2X1 U1819 ( .A(ram[862]), .B(n12982), .Y(n976) );
  OAI21X1 U1820 ( .A(n13056), .B(n12982), .C(n977), .Y(n5300) );
  NAND2X1 U1821 ( .A(ram[863]), .B(n12982), .Y(n977) );
  OAI21X1 U1823 ( .A(n13071), .B(n12981), .C(n979), .Y(n5301) );
  NAND2X1 U1824 ( .A(ram[864]), .B(n12981), .Y(n979) );
  OAI21X1 U1825 ( .A(n13070), .B(n12981), .C(n980), .Y(n5302) );
  NAND2X1 U1826 ( .A(ram[865]), .B(n12981), .Y(n980) );
  OAI21X1 U1827 ( .A(n13069), .B(n12981), .C(n981), .Y(n5303) );
  NAND2X1 U1828 ( .A(ram[866]), .B(n12981), .Y(n981) );
  OAI21X1 U1829 ( .A(n13068), .B(n12981), .C(n982), .Y(n5304) );
  NAND2X1 U1830 ( .A(ram[867]), .B(n12981), .Y(n982) );
  OAI21X1 U1831 ( .A(n13067), .B(n12981), .C(n983), .Y(n5305) );
  NAND2X1 U1832 ( .A(ram[868]), .B(n12981), .Y(n983) );
  OAI21X1 U1833 ( .A(n13066), .B(n12981), .C(n984), .Y(n5306) );
  NAND2X1 U1834 ( .A(ram[869]), .B(n12981), .Y(n984) );
  OAI21X1 U1835 ( .A(n13065), .B(n12981), .C(n985), .Y(n5307) );
  NAND2X1 U1836 ( .A(ram[870]), .B(n12981), .Y(n985) );
  OAI21X1 U1837 ( .A(n13064), .B(n12981), .C(n986), .Y(n5308) );
  NAND2X1 U1838 ( .A(ram[871]), .B(n12981), .Y(n986) );
  OAI21X1 U1839 ( .A(n13063), .B(n12981), .C(n987), .Y(n5309) );
  NAND2X1 U1840 ( .A(ram[872]), .B(n12981), .Y(n987) );
  OAI21X1 U1841 ( .A(n13062), .B(n12981), .C(n988), .Y(n5310) );
  NAND2X1 U1842 ( .A(ram[873]), .B(n12981), .Y(n988) );
  OAI21X1 U1843 ( .A(n13061), .B(n12981), .C(n989), .Y(n5311) );
  NAND2X1 U1844 ( .A(ram[874]), .B(n12981), .Y(n989) );
  OAI21X1 U1845 ( .A(n13060), .B(n12981), .C(n990), .Y(n5312) );
  NAND2X1 U1846 ( .A(ram[875]), .B(n12981), .Y(n990) );
  OAI21X1 U1847 ( .A(n13059), .B(n12981), .C(n991), .Y(n5313) );
  NAND2X1 U1848 ( .A(ram[876]), .B(n12981), .Y(n991) );
  OAI21X1 U1849 ( .A(n13058), .B(n12981), .C(n992), .Y(n5314) );
  NAND2X1 U1850 ( .A(ram[877]), .B(n12981), .Y(n992) );
  OAI21X1 U1851 ( .A(n13057), .B(n12981), .C(n993), .Y(n5315) );
  NAND2X1 U1852 ( .A(ram[878]), .B(n12981), .Y(n993) );
  OAI21X1 U1853 ( .A(n13056), .B(n12981), .C(n994), .Y(n5316) );
  NAND2X1 U1854 ( .A(ram[879]), .B(n12981), .Y(n994) );
  OAI21X1 U1856 ( .A(n12774), .B(n12980), .C(n996), .Y(n5317) );
  NAND2X1 U1857 ( .A(ram[880]), .B(n12980), .Y(n996) );
  OAI21X1 U1858 ( .A(n12768), .B(n12980), .C(n997), .Y(n5318) );
  NAND2X1 U1859 ( .A(ram[881]), .B(n12980), .Y(n997) );
  OAI21X1 U1860 ( .A(n13069), .B(n12980), .C(n998), .Y(n5319) );
  NAND2X1 U1861 ( .A(ram[882]), .B(n12980), .Y(n998) );
  OAI21X1 U1862 ( .A(n13068), .B(n12980), .C(n999), .Y(n5320) );
  NAND2X1 U1863 ( .A(ram[883]), .B(n12980), .Y(n999) );
  OAI21X1 U1864 ( .A(n13067), .B(n12980), .C(n1000), .Y(n5321) );
  NAND2X1 U1865 ( .A(ram[884]), .B(n12980), .Y(n1000) );
  OAI21X1 U1866 ( .A(n13066), .B(n12980), .C(n1001), .Y(n5322) );
  NAND2X1 U1867 ( .A(ram[885]), .B(n12980), .Y(n1001) );
  OAI21X1 U1868 ( .A(n13065), .B(n12980), .C(n1002), .Y(n5323) );
  NAND2X1 U1869 ( .A(ram[886]), .B(n12980), .Y(n1002) );
  OAI21X1 U1870 ( .A(n13064), .B(n12980), .C(n1003), .Y(n5324) );
  NAND2X1 U1871 ( .A(ram[887]), .B(n12980), .Y(n1003) );
  OAI21X1 U1872 ( .A(n13063), .B(n12980), .C(n1004), .Y(n5325) );
  NAND2X1 U1873 ( .A(ram[888]), .B(n12980), .Y(n1004) );
  OAI21X1 U1874 ( .A(n13062), .B(n12980), .C(n1005), .Y(n5326) );
  NAND2X1 U1875 ( .A(ram[889]), .B(n12980), .Y(n1005) );
  OAI21X1 U1876 ( .A(n13061), .B(n12980), .C(n1006), .Y(n5327) );
  NAND2X1 U1877 ( .A(ram[890]), .B(n12980), .Y(n1006) );
  OAI21X1 U1878 ( .A(n13060), .B(n12980), .C(n1007), .Y(n5328) );
  NAND2X1 U1879 ( .A(ram[891]), .B(n12980), .Y(n1007) );
  OAI21X1 U1880 ( .A(n13059), .B(n12980), .C(n1008), .Y(n5329) );
  NAND2X1 U1881 ( .A(ram[892]), .B(n12980), .Y(n1008) );
  OAI21X1 U1882 ( .A(n13058), .B(n12980), .C(n1009), .Y(n5330) );
  NAND2X1 U1883 ( .A(ram[893]), .B(n12980), .Y(n1009) );
  OAI21X1 U1884 ( .A(n12690), .B(n12980), .C(n1010), .Y(n5331) );
  NAND2X1 U1885 ( .A(ram[894]), .B(n12980), .Y(n1010) );
  OAI21X1 U1886 ( .A(n12684), .B(n12980), .C(n1011), .Y(n5332) );
  NAND2X1 U1887 ( .A(ram[895]), .B(n12980), .Y(n1011) );
  OAI21X1 U1889 ( .A(n12774), .B(n12979), .C(n1013), .Y(n5333) );
  NAND2X1 U1890 ( .A(ram[896]), .B(n12979), .Y(n1013) );
  OAI21X1 U1891 ( .A(n12768), .B(n12979), .C(n1014), .Y(n5334) );
  NAND2X1 U1892 ( .A(ram[897]), .B(n12979), .Y(n1014) );
  OAI21X1 U1893 ( .A(n13069), .B(n12979), .C(n1015), .Y(n5335) );
  NAND2X1 U1894 ( .A(ram[898]), .B(n12979), .Y(n1015) );
  OAI21X1 U1895 ( .A(n13068), .B(n12979), .C(n1016), .Y(n5336) );
  NAND2X1 U1896 ( .A(ram[899]), .B(n12979), .Y(n1016) );
  OAI21X1 U1897 ( .A(n13067), .B(n12979), .C(n1017), .Y(n5337) );
  NAND2X1 U1898 ( .A(ram[900]), .B(n12979), .Y(n1017) );
  OAI21X1 U1899 ( .A(n13066), .B(n12979), .C(n1018), .Y(n5338) );
  NAND2X1 U1900 ( .A(ram[901]), .B(n12979), .Y(n1018) );
  OAI21X1 U1901 ( .A(n13065), .B(n12979), .C(n1019), .Y(n5339) );
  NAND2X1 U1902 ( .A(ram[902]), .B(n12979), .Y(n1019) );
  OAI21X1 U1903 ( .A(n13064), .B(n12979), .C(n1020), .Y(n5340) );
  NAND2X1 U1904 ( .A(ram[903]), .B(n12979), .Y(n1020) );
  OAI21X1 U1905 ( .A(n13063), .B(n12979), .C(n1021), .Y(n5341) );
  NAND2X1 U1906 ( .A(ram[904]), .B(n12979), .Y(n1021) );
  OAI21X1 U1907 ( .A(n13062), .B(n12979), .C(n1022), .Y(n5342) );
  NAND2X1 U1908 ( .A(ram[905]), .B(n12979), .Y(n1022) );
  OAI21X1 U1909 ( .A(n13061), .B(n12979), .C(n1023), .Y(n5343) );
  NAND2X1 U1910 ( .A(ram[906]), .B(n12979), .Y(n1023) );
  OAI21X1 U1911 ( .A(n13060), .B(n12979), .C(n1024), .Y(n5344) );
  NAND2X1 U1912 ( .A(ram[907]), .B(n12979), .Y(n1024) );
  OAI21X1 U1913 ( .A(n13059), .B(n12979), .C(n1025), .Y(n5345) );
  NAND2X1 U1914 ( .A(ram[908]), .B(n12979), .Y(n1025) );
  OAI21X1 U1915 ( .A(n13058), .B(n12979), .C(n1026), .Y(n5346) );
  NAND2X1 U1916 ( .A(ram[909]), .B(n12979), .Y(n1026) );
  OAI21X1 U1917 ( .A(n12690), .B(n12979), .C(n1027), .Y(n5347) );
  NAND2X1 U1918 ( .A(ram[910]), .B(n12979), .Y(n1027) );
  OAI21X1 U1919 ( .A(n12684), .B(n12979), .C(n1028), .Y(n5348) );
  NAND2X1 U1920 ( .A(ram[911]), .B(n12979), .Y(n1028) );
  OAI21X1 U1922 ( .A(n12775), .B(n12978), .C(n1030), .Y(n5349) );
  NAND2X1 U1923 ( .A(ram[912]), .B(n12978), .Y(n1030) );
  OAI21X1 U1924 ( .A(n12769), .B(n12978), .C(n1031), .Y(n5350) );
  NAND2X1 U1925 ( .A(ram[913]), .B(n12978), .Y(n1031) );
  OAI21X1 U1926 ( .A(n13069), .B(n12978), .C(n1032), .Y(n5351) );
  NAND2X1 U1927 ( .A(ram[914]), .B(n12978), .Y(n1032) );
  OAI21X1 U1928 ( .A(n13068), .B(n12978), .C(n1033), .Y(n5352) );
  NAND2X1 U1929 ( .A(ram[915]), .B(n12978), .Y(n1033) );
  OAI21X1 U1930 ( .A(n13067), .B(n12978), .C(n1034), .Y(n5353) );
  NAND2X1 U1931 ( .A(ram[916]), .B(n12978), .Y(n1034) );
  OAI21X1 U1932 ( .A(n13066), .B(n12978), .C(n1035), .Y(n5354) );
  NAND2X1 U1933 ( .A(ram[917]), .B(n12978), .Y(n1035) );
  OAI21X1 U1934 ( .A(n13065), .B(n12978), .C(n1036), .Y(n5355) );
  NAND2X1 U1935 ( .A(ram[918]), .B(n12978), .Y(n1036) );
  OAI21X1 U1936 ( .A(n13064), .B(n12978), .C(n1037), .Y(n5356) );
  NAND2X1 U1937 ( .A(ram[919]), .B(n12978), .Y(n1037) );
  OAI21X1 U1938 ( .A(n13063), .B(n12978), .C(n1038), .Y(n5357) );
  NAND2X1 U1939 ( .A(ram[920]), .B(n12978), .Y(n1038) );
  OAI21X1 U1940 ( .A(n13062), .B(n12978), .C(n1039), .Y(n5358) );
  NAND2X1 U1941 ( .A(ram[921]), .B(n12978), .Y(n1039) );
  OAI21X1 U1942 ( .A(n13061), .B(n12978), .C(n1040), .Y(n5359) );
  NAND2X1 U1943 ( .A(ram[922]), .B(n12978), .Y(n1040) );
  OAI21X1 U1944 ( .A(n13060), .B(n12978), .C(n1041), .Y(n5360) );
  NAND2X1 U1945 ( .A(ram[923]), .B(n12978), .Y(n1041) );
  OAI21X1 U1946 ( .A(n13059), .B(n12978), .C(n1042), .Y(n5361) );
  NAND2X1 U1947 ( .A(ram[924]), .B(n12978), .Y(n1042) );
  OAI21X1 U1948 ( .A(n13058), .B(n12978), .C(n1043), .Y(n5362) );
  NAND2X1 U1949 ( .A(ram[925]), .B(n12978), .Y(n1043) );
  OAI21X1 U1950 ( .A(n12691), .B(n12978), .C(n1044), .Y(n5363) );
  NAND2X1 U1951 ( .A(ram[926]), .B(n12978), .Y(n1044) );
  OAI21X1 U1952 ( .A(n12685), .B(n12978), .C(n1045), .Y(n5364) );
  NAND2X1 U1953 ( .A(ram[927]), .B(n12978), .Y(n1045) );
  OAI21X1 U1955 ( .A(n12775), .B(n12977), .C(n1047), .Y(n5365) );
  NAND2X1 U1956 ( .A(ram[928]), .B(n12977), .Y(n1047) );
  OAI21X1 U1957 ( .A(n12769), .B(n12977), .C(n1048), .Y(n5366) );
  NAND2X1 U1958 ( .A(ram[929]), .B(n12977), .Y(n1048) );
  OAI21X1 U1959 ( .A(n12762), .B(n12977), .C(n1049), .Y(n5367) );
  NAND2X1 U1960 ( .A(ram[930]), .B(n12977), .Y(n1049) );
  OAI21X1 U1961 ( .A(n12756), .B(n12977), .C(n1050), .Y(n5368) );
  NAND2X1 U1962 ( .A(ram[931]), .B(n12977), .Y(n1050) );
  OAI21X1 U1963 ( .A(n12750), .B(n12977), .C(n1051), .Y(n5369) );
  NAND2X1 U1964 ( .A(ram[932]), .B(n12977), .Y(n1051) );
  OAI21X1 U1965 ( .A(n12744), .B(n12977), .C(n1052), .Y(n5370) );
  NAND2X1 U1966 ( .A(ram[933]), .B(n12977), .Y(n1052) );
  OAI21X1 U1967 ( .A(n12738), .B(n12977), .C(n1053), .Y(n5371) );
  NAND2X1 U1968 ( .A(ram[934]), .B(n12977), .Y(n1053) );
  OAI21X1 U1969 ( .A(n12732), .B(n12977), .C(n1054), .Y(n5372) );
  NAND2X1 U1970 ( .A(ram[935]), .B(n12977), .Y(n1054) );
  OAI21X1 U1971 ( .A(n12726), .B(n12977), .C(n1055), .Y(n5373) );
  NAND2X1 U1972 ( .A(ram[936]), .B(n12977), .Y(n1055) );
  OAI21X1 U1973 ( .A(n12720), .B(n12977), .C(n1056), .Y(n5374) );
  NAND2X1 U1974 ( .A(ram[937]), .B(n12977), .Y(n1056) );
  OAI21X1 U1975 ( .A(n12714), .B(n12977), .C(n1057), .Y(n5375) );
  NAND2X1 U1976 ( .A(ram[938]), .B(n12977), .Y(n1057) );
  OAI21X1 U1977 ( .A(n12708), .B(n12977), .C(n1058), .Y(n5376) );
  NAND2X1 U1978 ( .A(ram[939]), .B(n12977), .Y(n1058) );
  OAI21X1 U1979 ( .A(n12702), .B(n12977), .C(n1059), .Y(n5377) );
  NAND2X1 U1980 ( .A(ram[940]), .B(n12977), .Y(n1059) );
  OAI21X1 U1981 ( .A(n12696), .B(n12977), .C(n1060), .Y(n5378) );
  NAND2X1 U1982 ( .A(ram[941]), .B(n12977), .Y(n1060) );
  OAI21X1 U1983 ( .A(n12691), .B(n12977), .C(n1061), .Y(n5379) );
  NAND2X1 U1984 ( .A(ram[942]), .B(n12977), .Y(n1061) );
  OAI21X1 U1985 ( .A(n12685), .B(n12977), .C(n1062), .Y(n5380) );
  NAND2X1 U1986 ( .A(ram[943]), .B(n12977), .Y(n1062) );
  OAI21X1 U1988 ( .A(n12774), .B(n12976), .C(n1064), .Y(n5381) );
  NAND2X1 U1989 ( .A(ram[944]), .B(n12976), .Y(n1064) );
  OAI21X1 U1990 ( .A(n12768), .B(n12976), .C(n1065), .Y(n5382) );
  NAND2X1 U1991 ( .A(ram[945]), .B(n12976), .Y(n1065) );
  OAI21X1 U1992 ( .A(n12764), .B(n12976), .C(n1066), .Y(n5383) );
  NAND2X1 U1993 ( .A(ram[946]), .B(n12976), .Y(n1066) );
  OAI21X1 U1994 ( .A(n12758), .B(n12976), .C(n1067), .Y(n5384) );
  NAND2X1 U1995 ( .A(ram[947]), .B(n12976), .Y(n1067) );
  OAI21X1 U1996 ( .A(n12752), .B(n12976), .C(n1068), .Y(n5385) );
  NAND2X1 U1997 ( .A(ram[948]), .B(n12976), .Y(n1068) );
  OAI21X1 U1998 ( .A(n12746), .B(n12976), .C(n1069), .Y(n5386) );
  NAND2X1 U1999 ( .A(ram[949]), .B(n12976), .Y(n1069) );
  OAI21X1 U2000 ( .A(n12740), .B(n12976), .C(n1070), .Y(n5387) );
  NAND2X1 U2001 ( .A(ram[950]), .B(n12976), .Y(n1070) );
  OAI21X1 U2002 ( .A(n12734), .B(n12976), .C(n1071), .Y(n5388) );
  NAND2X1 U2003 ( .A(ram[951]), .B(n12976), .Y(n1071) );
  OAI21X1 U2004 ( .A(n12728), .B(n12976), .C(n1072), .Y(n5389) );
  NAND2X1 U2005 ( .A(ram[952]), .B(n12976), .Y(n1072) );
  OAI21X1 U2006 ( .A(n12722), .B(n12976), .C(n1073), .Y(n5390) );
  NAND2X1 U2007 ( .A(ram[953]), .B(n12976), .Y(n1073) );
  OAI21X1 U2008 ( .A(n12716), .B(n12976), .C(n1074), .Y(n5391) );
  NAND2X1 U2009 ( .A(ram[954]), .B(n12976), .Y(n1074) );
  OAI21X1 U2010 ( .A(n12710), .B(n12976), .C(n1075), .Y(n5392) );
  NAND2X1 U2011 ( .A(ram[955]), .B(n12976), .Y(n1075) );
  OAI21X1 U2012 ( .A(n12704), .B(n12976), .C(n1076), .Y(n5393) );
  NAND2X1 U2013 ( .A(ram[956]), .B(n12976), .Y(n1076) );
  OAI21X1 U2014 ( .A(n12698), .B(n12976), .C(n1077), .Y(n5394) );
  NAND2X1 U2015 ( .A(ram[957]), .B(n12976), .Y(n1077) );
  OAI21X1 U2016 ( .A(n12690), .B(n12976), .C(n1078), .Y(n5395) );
  NAND2X1 U2017 ( .A(ram[958]), .B(n12976), .Y(n1078) );
  OAI21X1 U2018 ( .A(n12684), .B(n12976), .C(n1079), .Y(n5396) );
  NAND2X1 U2019 ( .A(ram[959]), .B(n12976), .Y(n1079) );
  OAI21X1 U2021 ( .A(n13071), .B(n12975), .C(n1081), .Y(n5397) );
  NAND2X1 U2022 ( .A(ram[960]), .B(n12975), .Y(n1081) );
  OAI21X1 U2023 ( .A(n13070), .B(n12975), .C(n1082), .Y(n5398) );
  NAND2X1 U2024 ( .A(ram[961]), .B(n12975), .Y(n1082) );
  OAI21X1 U2025 ( .A(n12763), .B(n12975), .C(n1083), .Y(n5399) );
  NAND2X1 U2026 ( .A(ram[962]), .B(n12975), .Y(n1083) );
  OAI21X1 U2027 ( .A(n12757), .B(n12975), .C(n1084), .Y(n5400) );
  NAND2X1 U2028 ( .A(ram[963]), .B(n12975), .Y(n1084) );
  OAI21X1 U2029 ( .A(n12751), .B(n12975), .C(n1085), .Y(n5401) );
  NAND2X1 U2030 ( .A(ram[964]), .B(n12975), .Y(n1085) );
  OAI21X1 U2031 ( .A(n12745), .B(n12975), .C(n1086), .Y(n5402) );
  NAND2X1 U2032 ( .A(ram[965]), .B(n12975), .Y(n1086) );
  OAI21X1 U2033 ( .A(n12739), .B(n12975), .C(n1087), .Y(n5403) );
  NAND2X1 U2034 ( .A(ram[966]), .B(n12975), .Y(n1087) );
  OAI21X1 U2035 ( .A(n12733), .B(n12975), .C(n1088), .Y(n5404) );
  NAND2X1 U2036 ( .A(ram[967]), .B(n12975), .Y(n1088) );
  OAI21X1 U2037 ( .A(n12727), .B(n12975), .C(n1089), .Y(n5405) );
  NAND2X1 U2038 ( .A(ram[968]), .B(n12975), .Y(n1089) );
  OAI21X1 U2039 ( .A(n12721), .B(n12975), .C(n1090), .Y(n5406) );
  NAND2X1 U2040 ( .A(ram[969]), .B(n12975), .Y(n1090) );
  OAI21X1 U2041 ( .A(n12715), .B(n12975), .C(n1091), .Y(n5407) );
  NAND2X1 U2042 ( .A(ram[970]), .B(n12975), .Y(n1091) );
  OAI21X1 U2043 ( .A(n12709), .B(n12975), .C(n1092), .Y(n5408) );
  NAND2X1 U2044 ( .A(ram[971]), .B(n12975), .Y(n1092) );
  OAI21X1 U2045 ( .A(n12703), .B(n12975), .C(n1093), .Y(n5409) );
  NAND2X1 U2046 ( .A(ram[972]), .B(n12975), .Y(n1093) );
  OAI21X1 U2047 ( .A(n12697), .B(n12975), .C(n1094), .Y(n5410) );
  NAND2X1 U2048 ( .A(ram[973]), .B(n12975), .Y(n1094) );
  OAI21X1 U2049 ( .A(n13057), .B(n12975), .C(n1095), .Y(n5411) );
  NAND2X1 U2050 ( .A(ram[974]), .B(n12975), .Y(n1095) );
  OAI21X1 U2051 ( .A(n13056), .B(n12975), .C(n1096), .Y(n5412) );
  NAND2X1 U2052 ( .A(ram[975]), .B(n12975), .Y(n1096) );
  OAI21X1 U2054 ( .A(n13071), .B(n12974), .C(n1098), .Y(n5413) );
  NAND2X1 U2055 ( .A(ram[976]), .B(n12974), .Y(n1098) );
  OAI21X1 U2056 ( .A(n13070), .B(n12974), .C(n1099), .Y(n5414) );
  NAND2X1 U2057 ( .A(ram[977]), .B(n12974), .Y(n1099) );
  OAI21X1 U2058 ( .A(n12763), .B(n12974), .C(n1100), .Y(n5415) );
  NAND2X1 U2059 ( .A(ram[978]), .B(n12974), .Y(n1100) );
  OAI21X1 U2060 ( .A(n12757), .B(n12974), .C(n1101), .Y(n5416) );
  NAND2X1 U2061 ( .A(ram[979]), .B(n12974), .Y(n1101) );
  OAI21X1 U2062 ( .A(n12751), .B(n12974), .C(n1102), .Y(n5417) );
  NAND2X1 U2063 ( .A(ram[980]), .B(n12974), .Y(n1102) );
  OAI21X1 U2064 ( .A(n12745), .B(n12974), .C(n1103), .Y(n5418) );
  NAND2X1 U2065 ( .A(ram[981]), .B(n12974), .Y(n1103) );
  OAI21X1 U2066 ( .A(n12739), .B(n12974), .C(n1104), .Y(n5419) );
  NAND2X1 U2067 ( .A(ram[982]), .B(n12974), .Y(n1104) );
  OAI21X1 U2068 ( .A(n12733), .B(n12974), .C(n1105), .Y(n5420) );
  NAND2X1 U2069 ( .A(ram[983]), .B(n12974), .Y(n1105) );
  OAI21X1 U2070 ( .A(n12727), .B(n12974), .C(n1106), .Y(n5421) );
  NAND2X1 U2071 ( .A(ram[984]), .B(n12974), .Y(n1106) );
  OAI21X1 U2072 ( .A(n12721), .B(n12974), .C(n1107), .Y(n5422) );
  NAND2X1 U2073 ( .A(ram[985]), .B(n12974), .Y(n1107) );
  OAI21X1 U2074 ( .A(n12715), .B(n12974), .C(n1108), .Y(n5423) );
  NAND2X1 U2075 ( .A(ram[986]), .B(n12974), .Y(n1108) );
  OAI21X1 U2076 ( .A(n12709), .B(n12974), .C(n1109), .Y(n5424) );
  NAND2X1 U2077 ( .A(ram[987]), .B(n12974), .Y(n1109) );
  OAI21X1 U2078 ( .A(n12703), .B(n12974), .C(n1110), .Y(n5425) );
  NAND2X1 U2079 ( .A(ram[988]), .B(n12974), .Y(n1110) );
  OAI21X1 U2080 ( .A(n12697), .B(n12974), .C(n1111), .Y(n5426) );
  NAND2X1 U2081 ( .A(ram[989]), .B(n12974), .Y(n1111) );
  OAI21X1 U2082 ( .A(n13057), .B(n12974), .C(n1112), .Y(n5427) );
  NAND2X1 U2083 ( .A(ram[990]), .B(n12974), .Y(n1112) );
  OAI21X1 U2084 ( .A(n13056), .B(n12974), .C(n1113), .Y(n5428) );
  NAND2X1 U2085 ( .A(ram[991]), .B(n12974), .Y(n1113) );
  OAI21X1 U2087 ( .A(n12775), .B(n12973), .C(n1115), .Y(n5429) );
  NAND2X1 U2088 ( .A(ram[992]), .B(n12973), .Y(n1115) );
  OAI21X1 U2089 ( .A(n12769), .B(n12973), .C(n1116), .Y(n5430) );
  NAND2X1 U2090 ( .A(ram[993]), .B(n12973), .Y(n1116) );
  OAI21X1 U2091 ( .A(n13069), .B(n12973), .C(n1117), .Y(n5431) );
  NAND2X1 U2092 ( .A(ram[994]), .B(n12973), .Y(n1117) );
  OAI21X1 U2093 ( .A(n13068), .B(n12973), .C(n1118), .Y(n5432) );
  NAND2X1 U2094 ( .A(ram[995]), .B(n12973), .Y(n1118) );
  OAI21X1 U2095 ( .A(n13067), .B(n12973), .C(n1119), .Y(n5433) );
  NAND2X1 U2096 ( .A(ram[996]), .B(n12973), .Y(n1119) );
  OAI21X1 U2097 ( .A(n13066), .B(n12973), .C(n1120), .Y(n5434) );
  NAND2X1 U2098 ( .A(ram[997]), .B(n12973), .Y(n1120) );
  OAI21X1 U2099 ( .A(n13065), .B(n12973), .C(n1121), .Y(n5435) );
  NAND2X1 U2100 ( .A(ram[998]), .B(n12973), .Y(n1121) );
  OAI21X1 U2101 ( .A(n13064), .B(n12973), .C(n1122), .Y(n5436) );
  NAND2X1 U2102 ( .A(ram[999]), .B(n12973), .Y(n1122) );
  OAI21X1 U2103 ( .A(n13063), .B(n12973), .C(n1123), .Y(n5437) );
  NAND2X1 U2104 ( .A(ram[1000]), .B(n12973), .Y(n1123) );
  OAI21X1 U2105 ( .A(n13062), .B(n12973), .C(n1124), .Y(n5438) );
  NAND2X1 U2106 ( .A(ram[1001]), .B(n12973), .Y(n1124) );
  OAI21X1 U2107 ( .A(n13061), .B(n12973), .C(n1125), .Y(n5439) );
  NAND2X1 U2108 ( .A(ram[1002]), .B(n12973), .Y(n1125) );
  OAI21X1 U2109 ( .A(n13060), .B(n12973), .C(n1126), .Y(n5440) );
  NAND2X1 U2110 ( .A(ram[1003]), .B(n12973), .Y(n1126) );
  OAI21X1 U2111 ( .A(n13059), .B(n12973), .C(n1127), .Y(n5441) );
  NAND2X1 U2112 ( .A(ram[1004]), .B(n12973), .Y(n1127) );
  OAI21X1 U2113 ( .A(n13058), .B(n12973), .C(n1128), .Y(n5442) );
  NAND2X1 U2114 ( .A(ram[1005]), .B(n12973), .Y(n1128) );
  OAI21X1 U2115 ( .A(n12691), .B(n12973), .C(n1129), .Y(n5443) );
  NAND2X1 U2116 ( .A(ram[1006]), .B(n12973), .Y(n1129) );
  OAI21X1 U2117 ( .A(n12685), .B(n12973), .C(n1130), .Y(n5444) );
  NAND2X1 U2118 ( .A(ram[1007]), .B(n12973), .Y(n1130) );
  OAI21X1 U2120 ( .A(n12779), .B(n12972), .C(n1132), .Y(n5445) );
  NAND2X1 U2121 ( .A(ram[1008]), .B(n12972), .Y(n1132) );
  OAI21X1 U2122 ( .A(n12773), .B(n12972), .C(n1133), .Y(n5446) );
  NAND2X1 U2123 ( .A(ram[1009]), .B(n12972), .Y(n1133) );
  OAI21X1 U2124 ( .A(n12763), .B(n12972), .C(n1134), .Y(n5447) );
  NAND2X1 U2125 ( .A(ram[1010]), .B(n12972), .Y(n1134) );
  OAI21X1 U2126 ( .A(n12757), .B(n12972), .C(n1135), .Y(n5448) );
  NAND2X1 U2127 ( .A(ram[1011]), .B(n12972), .Y(n1135) );
  OAI21X1 U2128 ( .A(n12751), .B(n12972), .C(n1136), .Y(n5449) );
  NAND2X1 U2129 ( .A(ram[1012]), .B(n12972), .Y(n1136) );
  OAI21X1 U2130 ( .A(n12745), .B(n12972), .C(n1137), .Y(n5450) );
  NAND2X1 U2131 ( .A(ram[1013]), .B(n12972), .Y(n1137) );
  OAI21X1 U2132 ( .A(n12739), .B(n12972), .C(n1138), .Y(n5451) );
  NAND2X1 U2133 ( .A(ram[1014]), .B(n12972), .Y(n1138) );
  OAI21X1 U2134 ( .A(n12733), .B(n12972), .C(n1139), .Y(n5452) );
  NAND2X1 U2135 ( .A(ram[1015]), .B(n12972), .Y(n1139) );
  OAI21X1 U2136 ( .A(n12727), .B(n12972), .C(n1140), .Y(n5453) );
  NAND2X1 U2137 ( .A(ram[1016]), .B(n12972), .Y(n1140) );
  OAI21X1 U2138 ( .A(n12721), .B(n12972), .C(n1141), .Y(n5454) );
  NAND2X1 U2139 ( .A(ram[1017]), .B(n12972), .Y(n1141) );
  OAI21X1 U2140 ( .A(n12715), .B(n12972), .C(n1142), .Y(n5455) );
  NAND2X1 U2141 ( .A(ram[1018]), .B(n12972), .Y(n1142) );
  OAI21X1 U2142 ( .A(n12709), .B(n12972), .C(n1143), .Y(n5456) );
  NAND2X1 U2143 ( .A(ram[1019]), .B(n12972), .Y(n1143) );
  OAI21X1 U2144 ( .A(n12703), .B(n12972), .C(n1144), .Y(n5457) );
  NAND2X1 U2145 ( .A(ram[1020]), .B(n12972), .Y(n1144) );
  OAI21X1 U2146 ( .A(n12697), .B(n12972), .C(n1145), .Y(n5458) );
  NAND2X1 U2147 ( .A(ram[1021]), .B(n12972), .Y(n1145) );
  OAI21X1 U2148 ( .A(n12695), .B(n12972), .C(n1146), .Y(n5459) );
  NAND2X1 U2149 ( .A(ram[1022]), .B(n12972), .Y(n1146) );
  OAI21X1 U2150 ( .A(n12689), .B(n12972), .C(n1147), .Y(n5460) );
  NAND2X1 U2151 ( .A(ram[1023]), .B(n12972), .Y(n1147) );
  NAND3X1 U2153 ( .A(mem_write_en), .B(n326), .C(n1149), .Y(n1148) );
  NOR2X1 U2154 ( .A(mem_access_addr[6]), .B(mem_access_addr[7]), .Y(n326) );
  OAI21X1 U2155 ( .A(n13071), .B(n12971), .C(n1151), .Y(n5461) );
  NAND2X1 U2156 ( .A(ram[1024]), .B(n12971), .Y(n1151) );
  OAI21X1 U2157 ( .A(n13070), .B(n12971), .C(n1152), .Y(n5462) );
  NAND2X1 U2158 ( .A(ram[1025]), .B(n12971), .Y(n1152) );
  OAI21X1 U2159 ( .A(n13069), .B(n12971), .C(n1153), .Y(n5463) );
  NAND2X1 U2160 ( .A(ram[1026]), .B(n12971), .Y(n1153) );
  OAI21X1 U2161 ( .A(n13068), .B(n12971), .C(n1154), .Y(n5464) );
  NAND2X1 U2162 ( .A(ram[1027]), .B(n12971), .Y(n1154) );
  OAI21X1 U2163 ( .A(n13067), .B(n12971), .C(n1155), .Y(n5465) );
  NAND2X1 U2164 ( .A(ram[1028]), .B(n12971), .Y(n1155) );
  OAI21X1 U2165 ( .A(n13066), .B(n12971), .C(n1156), .Y(n5466) );
  NAND2X1 U2166 ( .A(ram[1029]), .B(n12971), .Y(n1156) );
  OAI21X1 U2167 ( .A(n13065), .B(n12971), .C(n1157), .Y(n5467) );
  NAND2X1 U2168 ( .A(ram[1030]), .B(n12971), .Y(n1157) );
  OAI21X1 U2169 ( .A(n13064), .B(n12971), .C(n1158), .Y(n5468) );
  NAND2X1 U2170 ( .A(ram[1031]), .B(n12971), .Y(n1158) );
  OAI21X1 U2171 ( .A(n13063), .B(n12971), .C(n1159), .Y(n5469) );
  NAND2X1 U2172 ( .A(ram[1032]), .B(n12971), .Y(n1159) );
  OAI21X1 U2173 ( .A(n13062), .B(n12971), .C(n1160), .Y(n5470) );
  NAND2X1 U2174 ( .A(ram[1033]), .B(n12971), .Y(n1160) );
  OAI21X1 U2175 ( .A(n13061), .B(n12971), .C(n1161), .Y(n5471) );
  NAND2X1 U2176 ( .A(ram[1034]), .B(n12971), .Y(n1161) );
  OAI21X1 U2177 ( .A(n13060), .B(n12971), .C(n1162), .Y(n5472) );
  NAND2X1 U2178 ( .A(ram[1035]), .B(n12971), .Y(n1162) );
  OAI21X1 U2179 ( .A(n13059), .B(n12971), .C(n1163), .Y(n5473) );
  NAND2X1 U2180 ( .A(ram[1036]), .B(n12971), .Y(n1163) );
  OAI21X1 U2181 ( .A(n13058), .B(n12971), .C(n1164), .Y(n5474) );
  NAND2X1 U2182 ( .A(ram[1037]), .B(n12971), .Y(n1164) );
  OAI21X1 U2183 ( .A(n13057), .B(n12971), .C(n1165), .Y(n5475) );
  NAND2X1 U2184 ( .A(ram[1038]), .B(n12971), .Y(n1165) );
  OAI21X1 U2185 ( .A(n13056), .B(n12971), .C(n1166), .Y(n5476) );
  NAND2X1 U2186 ( .A(ram[1039]), .B(n12971), .Y(n1166) );
  OAI21X1 U2188 ( .A(n13071), .B(n12970), .C(n1168), .Y(n5477) );
  NAND2X1 U2189 ( .A(ram[1040]), .B(n12970), .Y(n1168) );
  OAI21X1 U2190 ( .A(n13070), .B(n12970), .C(n1169), .Y(n5478) );
  NAND2X1 U2191 ( .A(ram[1041]), .B(n12970), .Y(n1169) );
  OAI21X1 U2192 ( .A(n13069), .B(n12970), .C(n1170), .Y(n5479) );
  NAND2X1 U2193 ( .A(ram[1042]), .B(n12970), .Y(n1170) );
  OAI21X1 U2194 ( .A(n13068), .B(n12970), .C(n1171), .Y(n5480) );
  NAND2X1 U2195 ( .A(ram[1043]), .B(n12970), .Y(n1171) );
  OAI21X1 U2196 ( .A(n13067), .B(n12970), .C(n1172), .Y(n5481) );
  NAND2X1 U2197 ( .A(ram[1044]), .B(n12970), .Y(n1172) );
  OAI21X1 U2198 ( .A(n13066), .B(n12970), .C(n1173), .Y(n5482) );
  NAND2X1 U2199 ( .A(ram[1045]), .B(n12970), .Y(n1173) );
  OAI21X1 U2200 ( .A(n13065), .B(n12970), .C(n1174), .Y(n5483) );
  NAND2X1 U2201 ( .A(ram[1046]), .B(n12970), .Y(n1174) );
  OAI21X1 U2202 ( .A(n13064), .B(n12970), .C(n1175), .Y(n5484) );
  NAND2X1 U2203 ( .A(ram[1047]), .B(n12970), .Y(n1175) );
  OAI21X1 U2204 ( .A(n13063), .B(n12970), .C(n1176), .Y(n5485) );
  NAND2X1 U2205 ( .A(ram[1048]), .B(n12970), .Y(n1176) );
  OAI21X1 U2206 ( .A(n13062), .B(n12970), .C(n1177), .Y(n5486) );
  NAND2X1 U2207 ( .A(ram[1049]), .B(n12970), .Y(n1177) );
  OAI21X1 U2208 ( .A(n13061), .B(n12970), .C(n1178), .Y(n5487) );
  NAND2X1 U2209 ( .A(ram[1050]), .B(n12970), .Y(n1178) );
  OAI21X1 U2210 ( .A(n13060), .B(n12970), .C(n1179), .Y(n5488) );
  NAND2X1 U2211 ( .A(ram[1051]), .B(n12970), .Y(n1179) );
  OAI21X1 U2212 ( .A(n13059), .B(n12970), .C(n1180), .Y(n5489) );
  NAND2X1 U2213 ( .A(ram[1052]), .B(n12970), .Y(n1180) );
  OAI21X1 U2214 ( .A(n13058), .B(n12970), .C(n1181), .Y(n5490) );
  NAND2X1 U2215 ( .A(ram[1053]), .B(n12970), .Y(n1181) );
  OAI21X1 U2216 ( .A(n13057), .B(n12970), .C(n1182), .Y(n5491) );
  NAND2X1 U2217 ( .A(ram[1054]), .B(n12970), .Y(n1182) );
  OAI21X1 U2218 ( .A(n13056), .B(n12970), .C(n1183), .Y(n5492) );
  NAND2X1 U2219 ( .A(ram[1055]), .B(n12970), .Y(n1183) );
  OAI21X1 U2221 ( .A(n13071), .B(n12969), .C(n1185), .Y(n5493) );
  NAND2X1 U2222 ( .A(ram[1056]), .B(n12969), .Y(n1185) );
  OAI21X1 U2223 ( .A(n13070), .B(n12969), .C(n1186), .Y(n5494) );
  NAND2X1 U2224 ( .A(ram[1057]), .B(n12969), .Y(n1186) );
  OAI21X1 U2225 ( .A(n13069), .B(n12969), .C(n1187), .Y(n5495) );
  NAND2X1 U2226 ( .A(ram[1058]), .B(n12969), .Y(n1187) );
  OAI21X1 U2227 ( .A(n13068), .B(n12969), .C(n1188), .Y(n5496) );
  NAND2X1 U2228 ( .A(ram[1059]), .B(n12969), .Y(n1188) );
  OAI21X1 U2229 ( .A(n13067), .B(n12969), .C(n1189), .Y(n5497) );
  NAND2X1 U2230 ( .A(ram[1060]), .B(n12969), .Y(n1189) );
  OAI21X1 U2231 ( .A(n13066), .B(n12969), .C(n1190), .Y(n5498) );
  NAND2X1 U2232 ( .A(ram[1061]), .B(n12969), .Y(n1190) );
  OAI21X1 U2233 ( .A(n13065), .B(n12969), .C(n1191), .Y(n5499) );
  NAND2X1 U2234 ( .A(ram[1062]), .B(n12969), .Y(n1191) );
  OAI21X1 U2235 ( .A(n13064), .B(n12969), .C(n1192), .Y(n5500) );
  NAND2X1 U2236 ( .A(ram[1063]), .B(n12969), .Y(n1192) );
  OAI21X1 U2237 ( .A(n13063), .B(n12969), .C(n1193), .Y(n5501) );
  NAND2X1 U2238 ( .A(ram[1064]), .B(n12969), .Y(n1193) );
  OAI21X1 U2239 ( .A(n13062), .B(n12969), .C(n1194), .Y(n5502) );
  NAND2X1 U2240 ( .A(ram[1065]), .B(n12969), .Y(n1194) );
  OAI21X1 U2241 ( .A(n13061), .B(n12969), .C(n1195), .Y(n5503) );
  NAND2X1 U2242 ( .A(ram[1066]), .B(n12969), .Y(n1195) );
  OAI21X1 U2243 ( .A(n13060), .B(n12969), .C(n1196), .Y(n5504) );
  NAND2X1 U2244 ( .A(ram[1067]), .B(n12969), .Y(n1196) );
  OAI21X1 U2245 ( .A(n13059), .B(n12969), .C(n1197), .Y(n5505) );
  NAND2X1 U2246 ( .A(ram[1068]), .B(n12969), .Y(n1197) );
  OAI21X1 U2247 ( .A(n13058), .B(n12969), .C(n1198), .Y(n5506) );
  NAND2X1 U2248 ( .A(ram[1069]), .B(n12969), .Y(n1198) );
  OAI21X1 U2249 ( .A(n13057), .B(n12969), .C(n1199), .Y(n5507) );
  NAND2X1 U2250 ( .A(ram[1070]), .B(n12969), .Y(n1199) );
  OAI21X1 U2251 ( .A(n13056), .B(n12969), .C(n1200), .Y(n5508) );
  NAND2X1 U2252 ( .A(ram[1071]), .B(n12969), .Y(n1200) );
  OAI21X1 U2254 ( .A(n12774), .B(n12968), .C(n1202), .Y(n5509) );
  NAND2X1 U2255 ( .A(ram[1072]), .B(n12968), .Y(n1202) );
  OAI21X1 U2256 ( .A(n12768), .B(n12968), .C(n1203), .Y(n5510) );
  NAND2X1 U2257 ( .A(ram[1073]), .B(n12968), .Y(n1203) );
  OAI21X1 U2258 ( .A(n12762), .B(n12968), .C(n1204), .Y(n5511) );
  NAND2X1 U2259 ( .A(ram[1074]), .B(n12968), .Y(n1204) );
  OAI21X1 U2260 ( .A(n12756), .B(n12968), .C(n1205), .Y(n5512) );
  NAND2X1 U2261 ( .A(ram[1075]), .B(n12968), .Y(n1205) );
  OAI21X1 U2262 ( .A(n12750), .B(n12968), .C(n1206), .Y(n5513) );
  NAND2X1 U2263 ( .A(ram[1076]), .B(n12968), .Y(n1206) );
  OAI21X1 U2264 ( .A(n12744), .B(n12968), .C(n1207), .Y(n5514) );
  NAND2X1 U2265 ( .A(ram[1077]), .B(n12968), .Y(n1207) );
  OAI21X1 U2266 ( .A(n12738), .B(n12968), .C(n1208), .Y(n5515) );
  NAND2X1 U2267 ( .A(ram[1078]), .B(n12968), .Y(n1208) );
  OAI21X1 U2268 ( .A(n12732), .B(n12968), .C(n1209), .Y(n5516) );
  NAND2X1 U2269 ( .A(ram[1079]), .B(n12968), .Y(n1209) );
  OAI21X1 U2270 ( .A(n12726), .B(n12968), .C(n1210), .Y(n5517) );
  NAND2X1 U2271 ( .A(ram[1080]), .B(n12968), .Y(n1210) );
  OAI21X1 U2272 ( .A(n12720), .B(n12968), .C(n1211), .Y(n5518) );
  NAND2X1 U2273 ( .A(ram[1081]), .B(n12968), .Y(n1211) );
  OAI21X1 U2274 ( .A(n12714), .B(n12968), .C(n1212), .Y(n5519) );
  NAND2X1 U2275 ( .A(ram[1082]), .B(n12968), .Y(n1212) );
  OAI21X1 U2276 ( .A(n12708), .B(n12968), .C(n1213), .Y(n5520) );
  NAND2X1 U2277 ( .A(ram[1083]), .B(n12968), .Y(n1213) );
  OAI21X1 U2278 ( .A(n12702), .B(n12968), .C(n1214), .Y(n5521) );
  NAND2X1 U2279 ( .A(ram[1084]), .B(n12968), .Y(n1214) );
  OAI21X1 U2280 ( .A(n12696), .B(n12968), .C(n1215), .Y(n5522) );
  NAND2X1 U2281 ( .A(ram[1085]), .B(n12968), .Y(n1215) );
  OAI21X1 U2282 ( .A(n12690), .B(n12968), .C(n1216), .Y(n5523) );
  NAND2X1 U2283 ( .A(ram[1086]), .B(n12968), .Y(n1216) );
  OAI21X1 U2284 ( .A(n12684), .B(n12968), .C(n1217), .Y(n5524) );
  NAND2X1 U2285 ( .A(ram[1087]), .B(n12968), .Y(n1217) );
  OAI21X1 U2287 ( .A(n12777), .B(n12967), .C(n1219), .Y(n5525) );
  NAND2X1 U2288 ( .A(ram[1088]), .B(n12967), .Y(n1219) );
  OAI21X1 U2289 ( .A(n12771), .B(n12967), .C(n1220), .Y(n5526) );
  NAND2X1 U2290 ( .A(ram[1089]), .B(n12967), .Y(n1220) );
  OAI21X1 U2291 ( .A(n12763), .B(n12967), .C(n1221), .Y(n5527) );
  NAND2X1 U2292 ( .A(ram[1090]), .B(n12967), .Y(n1221) );
  OAI21X1 U2293 ( .A(n12757), .B(n12967), .C(n1222), .Y(n5528) );
  NAND2X1 U2294 ( .A(ram[1091]), .B(n12967), .Y(n1222) );
  OAI21X1 U2295 ( .A(n12751), .B(n12967), .C(n1223), .Y(n5529) );
  NAND2X1 U2296 ( .A(ram[1092]), .B(n12967), .Y(n1223) );
  OAI21X1 U2297 ( .A(n12745), .B(n12967), .C(n1224), .Y(n5530) );
  NAND2X1 U2298 ( .A(ram[1093]), .B(n12967), .Y(n1224) );
  OAI21X1 U2299 ( .A(n12739), .B(n12967), .C(n1225), .Y(n5531) );
  NAND2X1 U2300 ( .A(ram[1094]), .B(n12967), .Y(n1225) );
  OAI21X1 U2301 ( .A(n12733), .B(n12967), .C(n1226), .Y(n5532) );
  NAND2X1 U2302 ( .A(ram[1095]), .B(n12967), .Y(n1226) );
  OAI21X1 U2303 ( .A(n12727), .B(n12967), .C(n1227), .Y(n5533) );
  NAND2X1 U2304 ( .A(ram[1096]), .B(n12967), .Y(n1227) );
  OAI21X1 U2305 ( .A(n12721), .B(n12967), .C(n1228), .Y(n5534) );
  NAND2X1 U2306 ( .A(ram[1097]), .B(n12967), .Y(n1228) );
  OAI21X1 U2307 ( .A(n12715), .B(n12967), .C(n1229), .Y(n5535) );
  NAND2X1 U2308 ( .A(ram[1098]), .B(n12967), .Y(n1229) );
  OAI21X1 U2309 ( .A(n12709), .B(n12967), .C(n1230), .Y(n5536) );
  NAND2X1 U2310 ( .A(ram[1099]), .B(n12967), .Y(n1230) );
  OAI21X1 U2311 ( .A(n12703), .B(n12967), .C(n1231), .Y(n5537) );
  NAND2X1 U2312 ( .A(ram[1100]), .B(n12967), .Y(n1231) );
  OAI21X1 U2313 ( .A(n12697), .B(n12967), .C(n1232), .Y(n5538) );
  NAND2X1 U2314 ( .A(ram[1101]), .B(n12967), .Y(n1232) );
  OAI21X1 U2315 ( .A(n12693), .B(n12967), .C(n1233), .Y(n5539) );
  NAND2X1 U2316 ( .A(ram[1102]), .B(n12967), .Y(n1233) );
  OAI21X1 U2317 ( .A(n12687), .B(n12967), .C(n1234), .Y(n5540) );
  NAND2X1 U2318 ( .A(ram[1103]), .B(n12967), .Y(n1234) );
  OAI21X1 U2320 ( .A(n12775), .B(n12966), .C(n1236), .Y(n5541) );
  NAND2X1 U2321 ( .A(ram[1104]), .B(n12966), .Y(n1236) );
  OAI21X1 U2322 ( .A(n12769), .B(n12966), .C(n1237), .Y(n5542) );
  NAND2X1 U2323 ( .A(ram[1105]), .B(n12966), .Y(n1237) );
  OAI21X1 U2324 ( .A(n12763), .B(n12966), .C(n1238), .Y(n5543) );
  NAND2X1 U2325 ( .A(ram[1106]), .B(n12966), .Y(n1238) );
  OAI21X1 U2326 ( .A(n12757), .B(n12966), .C(n1239), .Y(n5544) );
  NAND2X1 U2327 ( .A(ram[1107]), .B(n12966), .Y(n1239) );
  OAI21X1 U2328 ( .A(n12751), .B(n12966), .C(n1240), .Y(n5545) );
  NAND2X1 U2329 ( .A(ram[1108]), .B(n12966), .Y(n1240) );
  OAI21X1 U2330 ( .A(n12745), .B(n12966), .C(n1241), .Y(n5546) );
  NAND2X1 U2331 ( .A(ram[1109]), .B(n12966), .Y(n1241) );
  OAI21X1 U2332 ( .A(n12739), .B(n12966), .C(n1242), .Y(n5547) );
  NAND2X1 U2333 ( .A(ram[1110]), .B(n12966), .Y(n1242) );
  OAI21X1 U2334 ( .A(n12733), .B(n12966), .C(n1243), .Y(n5548) );
  NAND2X1 U2335 ( .A(ram[1111]), .B(n12966), .Y(n1243) );
  OAI21X1 U2336 ( .A(n12727), .B(n12966), .C(n1244), .Y(n5549) );
  NAND2X1 U2337 ( .A(ram[1112]), .B(n12966), .Y(n1244) );
  OAI21X1 U2338 ( .A(n12721), .B(n12966), .C(n1245), .Y(n5550) );
  NAND2X1 U2339 ( .A(ram[1113]), .B(n12966), .Y(n1245) );
  OAI21X1 U2340 ( .A(n12715), .B(n12966), .C(n1246), .Y(n5551) );
  NAND2X1 U2341 ( .A(ram[1114]), .B(n12966), .Y(n1246) );
  OAI21X1 U2342 ( .A(n12709), .B(n12966), .C(n1247), .Y(n5552) );
  NAND2X1 U2343 ( .A(ram[1115]), .B(n12966), .Y(n1247) );
  OAI21X1 U2344 ( .A(n12703), .B(n12966), .C(n1248), .Y(n5553) );
  NAND2X1 U2345 ( .A(ram[1116]), .B(n12966), .Y(n1248) );
  OAI21X1 U2346 ( .A(n12697), .B(n12966), .C(n1249), .Y(n5554) );
  NAND2X1 U2347 ( .A(ram[1117]), .B(n12966), .Y(n1249) );
  OAI21X1 U2348 ( .A(n12691), .B(n12966), .C(n1250), .Y(n5555) );
  NAND2X1 U2349 ( .A(ram[1118]), .B(n12966), .Y(n1250) );
  OAI21X1 U2350 ( .A(n12685), .B(n12966), .C(n1251), .Y(n5556) );
  NAND2X1 U2351 ( .A(ram[1119]), .B(n12966), .Y(n1251) );
  OAI21X1 U2353 ( .A(n12774), .B(n12965), .C(n1253), .Y(n5557) );
  NAND2X1 U2354 ( .A(ram[1120]), .B(n12965), .Y(n1253) );
  OAI21X1 U2355 ( .A(n12768), .B(n12965), .C(n1254), .Y(n5558) );
  NAND2X1 U2356 ( .A(ram[1121]), .B(n12965), .Y(n1254) );
  OAI21X1 U2357 ( .A(n12762), .B(n12965), .C(n1255), .Y(n5559) );
  NAND2X1 U2358 ( .A(ram[1122]), .B(n12965), .Y(n1255) );
  OAI21X1 U2359 ( .A(n12756), .B(n12965), .C(n1256), .Y(n5560) );
  NAND2X1 U2360 ( .A(ram[1123]), .B(n12965), .Y(n1256) );
  OAI21X1 U2361 ( .A(n12750), .B(n12965), .C(n1257), .Y(n5561) );
  NAND2X1 U2362 ( .A(ram[1124]), .B(n12965), .Y(n1257) );
  OAI21X1 U2363 ( .A(n12744), .B(n12965), .C(n1258), .Y(n5562) );
  NAND2X1 U2364 ( .A(ram[1125]), .B(n12965), .Y(n1258) );
  OAI21X1 U2365 ( .A(n12738), .B(n12965), .C(n1259), .Y(n5563) );
  NAND2X1 U2366 ( .A(ram[1126]), .B(n12965), .Y(n1259) );
  OAI21X1 U2367 ( .A(n12732), .B(n12965), .C(n1260), .Y(n5564) );
  NAND2X1 U2368 ( .A(ram[1127]), .B(n12965), .Y(n1260) );
  OAI21X1 U2369 ( .A(n12726), .B(n12965), .C(n1261), .Y(n5565) );
  NAND2X1 U2370 ( .A(ram[1128]), .B(n12965), .Y(n1261) );
  OAI21X1 U2371 ( .A(n12720), .B(n12965), .C(n1262), .Y(n5566) );
  NAND2X1 U2372 ( .A(ram[1129]), .B(n12965), .Y(n1262) );
  OAI21X1 U2373 ( .A(n12714), .B(n12965), .C(n1263), .Y(n5567) );
  NAND2X1 U2374 ( .A(ram[1130]), .B(n12965), .Y(n1263) );
  OAI21X1 U2375 ( .A(n12708), .B(n12965), .C(n1264), .Y(n5568) );
  NAND2X1 U2376 ( .A(ram[1131]), .B(n12965), .Y(n1264) );
  OAI21X1 U2377 ( .A(n12702), .B(n12965), .C(n1265), .Y(n5569) );
  NAND2X1 U2378 ( .A(ram[1132]), .B(n12965), .Y(n1265) );
  OAI21X1 U2379 ( .A(n12696), .B(n12965), .C(n1266), .Y(n5570) );
  NAND2X1 U2380 ( .A(ram[1133]), .B(n12965), .Y(n1266) );
  OAI21X1 U2381 ( .A(n12690), .B(n12965), .C(n1267), .Y(n5571) );
  NAND2X1 U2382 ( .A(ram[1134]), .B(n12965), .Y(n1267) );
  OAI21X1 U2383 ( .A(n12684), .B(n12965), .C(n1268), .Y(n5572) );
  NAND2X1 U2384 ( .A(ram[1135]), .B(n12965), .Y(n1268) );
  OAI21X1 U2386 ( .A(n12775), .B(n12964), .C(n1270), .Y(n5573) );
  NAND2X1 U2387 ( .A(ram[1136]), .B(n12964), .Y(n1270) );
  OAI21X1 U2388 ( .A(n12769), .B(n12964), .C(n1271), .Y(n5574) );
  NAND2X1 U2389 ( .A(ram[1137]), .B(n12964), .Y(n1271) );
  OAI21X1 U2390 ( .A(n12762), .B(n12964), .C(n1272), .Y(n5575) );
  NAND2X1 U2391 ( .A(ram[1138]), .B(n12964), .Y(n1272) );
  OAI21X1 U2392 ( .A(n12756), .B(n12964), .C(n1273), .Y(n5576) );
  NAND2X1 U2393 ( .A(ram[1139]), .B(n12964), .Y(n1273) );
  OAI21X1 U2394 ( .A(n12750), .B(n12964), .C(n1274), .Y(n5577) );
  NAND2X1 U2395 ( .A(ram[1140]), .B(n12964), .Y(n1274) );
  OAI21X1 U2396 ( .A(n12744), .B(n12964), .C(n1275), .Y(n5578) );
  NAND2X1 U2397 ( .A(ram[1141]), .B(n12964), .Y(n1275) );
  OAI21X1 U2398 ( .A(n12738), .B(n12964), .C(n1276), .Y(n5579) );
  NAND2X1 U2399 ( .A(ram[1142]), .B(n12964), .Y(n1276) );
  OAI21X1 U2400 ( .A(n12732), .B(n12964), .C(n1277), .Y(n5580) );
  NAND2X1 U2401 ( .A(ram[1143]), .B(n12964), .Y(n1277) );
  OAI21X1 U2402 ( .A(n12726), .B(n12964), .C(n1278), .Y(n5581) );
  NAND2X1 U2403 ( .A(ram[1144]), .B(n12964), .Y(n1278) );
  OAI21X1 U2404 ( .A(n12720), .B(n12964), .C(n1279), .Y(n5582) );
  NAND2X1 U2405 ( .A(ram[1145]), .B(n12964), .Y(n1279) );
  OAI21X1 U2406 ( .A(n12714), .B(n12964), .C(n1280), .Y(n5583) );
  NAND2X1 U2407 ( .A(ram[1146]), .B(n12964), .Y(n1280) );
  OAI21X1 U2408 ( .A(n12708), .B(n12964), .C(n1281), .Y(n5584) );
  NAND2X1 U2409 ( .A(ram[1147]), .B(n12964), .Y(n1281) );
  OAI21X1 U2410 ( .A(n12702), .B(n12964), .C(n1282), .Y(n5585) );
  NAND2X1 U2411 ( .A(ram[1148]), .B(n12964), .Y(n1282) );
  OAI21X1 U2412 ( .A(n12696), .B(n12964), .C(n1283), .Y(n5586) );
  NAND2X1 U2413 ( .A(ram[1149]), .B(n12964), .Y(n1283) );
  OAI21X1 U2414 ( .A(n12691), .B(n12964), .C(n1284), .Y(n5587) );
  NAND2X1 U2415 ( .A(ram[1150]), .B(n12964), .Y(n1284) );
  OAI21X1 U2416 ( .A(n12685), .B(n12964), .C(n1285), .Y(n5588) );
  NAND2X1 U2417 ( .A(ram[1151]), .B(n12964), .Y(n1285) );
  OAI21X1 U2419 ( .A(n12775), .B(n12963), .C(n1287), .Y(n5589) );
  NAND2X1 U2420 ( .A(ram[1152]), .B(n12963), .Y(n1287) );
  OAI21X1 U2421 ( .A(n12769), .B(n12963), .C(n1288), .Y(n5590) );
  NAND2X1 U2422 ( .A(ram[1153]), .B(n12963), .Y(n1288) );
  OAI21X1 U2423 ( .A(n12763), .B(n12963), .C(n1289), .Y(n5591) );
  NAND2X1 U2424 ( .A(ram[1154]), .B(n12963), .Y(n1289) );
  OAI21X1 U2425 ( .A(n12757), .B(n12963), .C(n1290), .Y(n5592) );
  NAND2X1 U2426 ( .A(ram[1155]), .B(n12963), .Y(n1290) );
  OAI21X1 U2427 ( .A(n12751), .B(n12963), .C(n1291), .Y(n5593) );
  NAND2X1 U2428 ( .A(ram[1156]), .B(n12963), .Y(n1291) );
  OAI21X1 U2429 ( .A(n12745), .B(n12963), .C(n1292), .Y(n5594) );
  NAND2X1 U2430 ( .A(ram[1157]), .B(n12963), .Y(n1292) );
  OAI21X1 U2431 ( .A(n12739), .B(n12963), .C(n1293), .Y(n5595) );
  NAND2X1 U2432 ( .A(ram[1158]), .B(n12963), .Y(n1293) );
  OAI21X1 U2433 ( .A(n12733), .B(n12963), .C(n1294), .Y(n5596) );
  NAND2X1 U2434 ( .A(ram[1159]), .B(n12963), .Y(n1294) );
  OAI21X1 U2435 ( .A(n12727), .B(n12963), .C(n1295), .Y(n5597) );
  NAND2X1 U2436 ( .A(ram[1160]), .B(n12963), .Y(n1295) );
  OAI21X1 U2437 ( .A(n12721), .B(n12963), .C(n1296), .Y(n5598) );
  NAND2X1 U2438 ( .A(ram[1161]), .B(n12963), .Y(n1296) );
  OAI21X1 U2439 ( .A(n12715), .B(n12963), .C(n1297), .Y(n5599) );
  NAND2X1 U2440 ( .A(ram[1162]), .B(n12963), .Y(n1297) );
  OAI21X1 U2441 ( .A(n12709), .B(n12963), .C(n1298), .Y(n5600) );
  NAND2X1 U2442 ( .A(ram[1163]), .B(n12963), .Y(n1298) );
  OAI21X1 U2443 ( .A(n12703), .B(n12963), .C(n1299), .Y(n5601) );
  NAND2X1 U2444 ( .A(ram[1164]), .B(n12963), .Y(n1299) );
  OAI21X1 U2445 ( .A(n12697), .B(n12963), .C(n1300), .Y(n5602) );
  NAND2X1 U2446 ( .A(ram[1165]), .B(n12963), .Y(n1300) );
  OAI21X1 U2447 ( .A(n12691), .B(n12963), .C(n1301), .Y(n5603) );
  NAND2X1 U2448 ( .A(ram[1166]), .B(n12963), .Y(n1301) );
  OAI21X1 U2449 ( .A(n12685), .B(n12963), .C(n1302), .Y(n5604) );
  NAND2X1 U2450 ( .A(ram[1167]), .B(n12963), .Y(n1302) );
  OAI21X1 U2452 ( .A(n13071), .B(n12962), .C(n1304), .Y(n5605) );
  NAND2X1 U2453 ( .A(ram[1168]), .B(n12962), .Y(n1304) );
  OAI21X1 U2454 ( .A(n13070), .B(n12962), .C(n1305), .Y(n5606) );
  NAND2X1 U2455 ( .A(ram[1169]), .B(n12962), .Y(n1305) );
  OAI21X1 U2456 ( .A(n13069), .B(n12962), .C(n1306), .Y(n5607) );
  NAND2X1 U2457 ( .A(ram[1170]), .B(n12962), .Y(n1306) );
  OAI21X1 U2458 ( .A(n13068), .B(n12962), .C(n1307), .Y(n5608) );
  NAND2X1 U2459 ( .A(ram[1171]), .B(n12962), .Y(n1307) );
  OAI21X1 U2460 ( .A(n13067), .B(n12962), .C(n1308), .Y(n5609) );
  NAND2X1 U2461 ( .A(ram[1172]), .B(n12962), .Y(n1308) );
  OAI21X1 U2462 ( .A(n13066), .B(n12962), .C(n1309), .Y(n5610) );
  NAND2X1 U2463 ( .A(ram[1173]), .B(n12962), .Y(n1309) );
  OAI21X1 U2464 ( .A(n13065), .B(n12962), .C(n1310), .Y(n5611) );
  NAND2X1 U2465 ( .A(ram[1174]), .B(n12962), .Y(n1310) );
  OAI21X1 U2466 ( .A(n13064), .B(n12962), .C(n1311), .Y(n5612) );
  NAND2X1 U2467 ( .A(ram[1175]), .B(n12962), .Y(n1311) );
  OAI21X1 U2468 ( .A(n13063), .B(n12962), .C(n1312), .Y(n5613) );
  NAND2X1 U2469 ( .A(ram[1176]), .B(n12962), .Y(n1312) );
  OAI21X1 U2470 ( .A(n13062), .B(n12962), .C(n1313), .Y(n5614) );
  NAND2X1 U2471 ( .A(ram[1177]), .B(n12962), .Y(n1313) );
  OAI21X1 U2472 ( .A(n13061), .B(n12962), .C(n1314), .Y(n5615) );
  NAND2X1 U2473 ( .A(ram[1178]), .B(n12962), .Y(n1314) );
  OAI21X1 U2474 ( .A(n13060), .B(n12962), .C(n1315), .Y(n5616) );
  NAND2X1 U2475 ( .A(ram[1179]), .B(n12962), .Y(n1315) );
  OAI21X1 U2476 ( .A(n13059), .B(n12962), .C(n1316), .Y(n5617) );
  NAND2X1 U2477 ( .A(ram[1180]), .B(n12962), .Y(n1316) );
  OAI21X1 U2478 ( .A(n13058), .B(n12962), .C(n1317), .Y(n5618) );
  NAND2X1 U2479 ( .A(ram[1181]), .B(n12962), .Y(n1317) );
  OAI21X1 U2480 ( .A(n13057), .B(n12962), .C(n1318), .Y(n5619) );
  NAND2X1 U2481 ( .A(ram[1182]), .B(n12962), .Y(n1318) );
  OAI21X1 U2482 ( .A(n13056), .B(n12962), .C(n1319), .Y(n5620) );
  NAND2X1 U2483 ( .A(ram[1183]), .B(n12962), .Y(n1319) );
  OAI21X1 U2485 ( .A(n12778), .B(n12961), .C(n1321), .Y(n5621) );
  NAND2X1 U2486 ( .A(ram[1184]), .B(n12961), .Y(n1321) );
  OAI21X1 U2487 ( .A(n12772), .B(n12961), .C(n1322), .Y(n5622) );
  NAND2X1 U2488 ( .A(ram[1185]), .B(n12961), .Y(n1322) );
  OAI21X1 U2489 ( .A(n12767), .B(n12961), .C(n1323), .Y(n5623) );
  NAND2X1 U2490 ( .A(ram[1186]), .B(n12961), .Y(n1323) );
  OAI21X1 U2491 ( .A(n12761), .B(n12961), .C(n1324), .Y(n5624) );
  NAND2X1 U2492 ( .A(ram[1187]), .B(n12961), .Y(n1324) );
  OAI21X1 U2493 ( .A(n12755), .B(n12961), .C(n1325), .Y(n5625) );
  NAND2X1 U2494 ( .A(ram[1188]), .B(n12961), .Y(n1325) );
  OAI21X1 U2495 ( .A(n12749), .B(n12961), .C(n1326), .Y(n5626) );
  NAND2X1 U2496 ( .A(ram[1189]), .B(n12961), .Y(n1326) );
  OAI21X1 U2497 ( .A(n12743), .B(n12961), .C(n1327), .Y(n5627) );
  NAND2X1 U2498 ( .A(ram[1190]), .B(n12961), .Y(n1327) );
  OAI21X1 U2499 ( .A(n12737), .B(n12961), .C(n1328), .Y(n5628) );
  NAND2X1 U2500 ( .A(ram[1191]), .B(n12961), .Y(n1328) );
  OAI21X1 U2501 ( .A(n12731), .B(n12961), .C(n1329), .Y(n5629) );
  NAND2X1 U2502 ( .A(ram[1192]), .B(n12961), .Y(n1329) );
  OAI21X1 U2503 ( .A(n12725), .B(n12961), .C(n1330), .Y(n5630) );
  NAND2X1 U2504 ( .A(ram[1193]), .B(n12961), .Y(n1330) );
  OAI21X1 U2505 ( .A(n12719), .B(n12961), .C(n1331), .Y(n5631) );
  NAND2X1 U2506 ( .A(ram[1194]), .B(n12961), .Y(n1331) );
  OAI21X1 U2507 ( .A(n12713), .B(n12961), .C(n1332), .Y(n5632) );
  NAND2X1 U2508 ( .A(ram[1195]), .B(n12961), .Y(n1332) );
  OAI21X1 U2509 ( .A(n12707), .B(n12961), .C(n1333), .Y(n5633) );
  NAND2X1 U2510 ( .A(ram[1196]), .B(n12961), .Y(n1333) );
  OAI21X1 U2511 ( .A(n12701), .B(n12961), .C(n1334), .Y(n5634) );
  NAND2X1 U2512 ( .A(ram[1197]), .B(n12961), .Y(n1334) );
  OAI21X1 U2513 ( .A(n12694), .B(n12961), .C(n1335), .Y(n5635) );
  NAND2X1 U2514 ( .A(ram[1198]), .B(n12961), .Y(n1335) );
  OAI21X1 U2515 ( .A(n12688), .B(n12961), .C(n1336), .Y(n5636) );
  NAND2X1 U2516 ( .A(ram[1199]), .B(n12961), .Y(n1336) );
  OAI21X1 U2518 ( .A(n12779), .B(n12960), .C(n1338), .Y(n5637) );
  NAND2X1 U2519 ( .A(ram[1200]), .B(n12960), .Y(n1338) );
  OAI21X1 U2520 ( .A(n12773), .B(n12960), .C(n1339), .Y(n5638) );
  NAND2X1 U2521 ( .A(ram[1201]), .B(n12960), .Y(n1339) );
  OAI21X1 U2522 ( .A(n12764), .B(n12960), .C(n1340), .Y(n5639) );
  NAND2X1 U2523 ( .A(ram[1202]), .B(n12960), .Y(n1340) );
  OAI21X1 U2524 ( .A(n12758), .B(n12960), .C(n1341), .Y(n5640) );
  NAND2X1 U2525 ( .A(ram[1203]), .B(n12960), .Y(n1341) );
  OAI21X1 U2526 ( .A(n12752), .B(n12960), .C(n1342), .Y(n5641) );
  NAND2X1 U2527 ( .A(ram[1204]), .B(n12960), .Y(n1342) );
  OAI21X1 U2528 ( .A(n12746), .B(n12960), .C(n1343), .Y(n5642) );
  NAND2X1 U2529 ( .A(ram[1205]), .B(n12960), .Y(n1343) );
  OAI21X1 U2530 ( .A(n12740), .B(n12960), .C(n1344), .Y(n5643) );
  NAND2X1 U2531 ( .A(ram[1206]), .B(n12960), .Y(n1344) );
  OAI21X1 U2532 ( .A(n12734), .B(n12960), .C(n1345), .Y(n5644) );
  NAND2X1 U2533 ( .A(ram[1207]), .B(n12960), .Y(n1345) );
  OAI21X1 U2534 ( .A(n12728), .B(n12960), .C(n1346), .Y(n5645) );
  NAND2X1 U2535 ( .A(ram[1208]), .B(n12960), .Y(n1346) );
  OAI21X1 U2536 ( .A(n12722), .B(n12960), .C(n1347), .Y(n5646) );
  NAND2X1 U2537 ( .A(ram[1209]), .B(n12960), .Y(n1347) );
  OAI21X1 U2538 ( .A(n12716), .B(n12960), .C(n1348), .Y(n5647) );
  NAND2X1 U2539 ( .A(ram[1210]), .B(n12960), .Y(n1348) );
  OAI21X1 U2540 ( .A(n12710), .B(n12960), .C(n1349), .Y(n5648) );
  NAND2X1 U2541 ( .A(ram[1211]), .B(n12960), .Y(n1349) );
  OAI21X1 U2542 ( .A(n12704), .B(n12960), .C(n1350), .Y(n5649) );
  NAND2X1 U2543 ( .A(ram[1212]), .B(n12960), .Y(n1350) );
  OAI21X1 U2544 ( .A(n12698), .B(n12960), .C(n1351), .Y(n5650) );
  NAND2X1 U2545 ( .A(ram[1213]), .B(n12960), .Y(n1351) );
  OAI21X1 U2546 ( .A(n12695), .B(n12960), .C(n1352), .Y(n5651) );
  NAND2X1 U2547 ( .A(ram[1214]), .B(n12960), .Y(n1352) );
  OAI21X1 U2548 ( .A(n12689), .B(n12960), .C(n1353), .Y(n5652) );
  NAND2X1 U2549 ( .A(ram[1215]), .B(n12960), .Y(n1353) );
  OAI21X1 U2551 ( .A(n12776), .B(n12959), .C(n1355), .Y(n5653) );
  NAND2X1 U2552 ( .A(ram[1216]), .B(n12959), .Y(n1355) );
  OAI21X1 U2553 ( .A(n12770), .B(n12959), .C(n1356), .Y(n5654) );
  NAND2X1 U2554 ( .A(ram[1217]), .B(n12959), .Y(n1356) );
  OAI21X1 U2555 ( .A(n12767), .B(n12959), .C(n1357), .Y(n5655) );
  NAND2X1 U2556 ( .A(ram[1218]), .B(n12959), .Y(n1357) );
  OAI21X1 U2557 ( .A(n12761), .B(n12959), .C(n1358), .Y(n5656) );
  NAND2X1 U2558 ( .A(ram[1219]), .B(n12959), .Y(n1358) );
  OAI21X1 U2559 ( .A(n12755), .B(n12959), .C(n1359), .Y(n5657) );
  NAND2X1 U2560 ( .A(ram[1220]), .B(n12959), .Y(n1359) );
  OAI21X1 U2561 ( .A(n12749), .B(n12959), .C(n1360), .Y(n5658) );
  NAND2X1 U2562 ( .A(ram[1221]), .B(n12959), .Y(n1360) );
  OAI21X1 U2563 ( .A(n12743), .B(n12959), .C(n1361), .Y(n5659) );
  NAND2X1 U2564 ( .A(ram[1222]), .B(n12959), .Y(n1361) );
  OAI21X1 U2565 ( .A(n12737), .B(n12959), .C(n1362), .Y(n5660) );
  NAND2X1 U2566 ( .A(ram[1223]), .B(n12959), .Y(n1362) );
  OAI21X1 U2567 ( .A(n12731), .B(n12959), .C(n1363), .Y(n5661) );
  NAND2X1 U2568 ( .A(ram[1224]), .B(n12959), .Y(n1363) );
  OAI21X1 U2569 ( .A(n12725), .B(n12959), .C(n1364), .Y(n5662) );
  NAND2X1 U2570 ( .A(ram[1225]), .B(n12959), .Y(n1364) );
  OAI21X1 U2571 ( .A(n12719), .B(n12959), .C(n1365), .Y(n5663) );
  NAND2X1 U2572 ( .A(ram[1226]), .B(n12959), .Y(n1365) );
  OAI21X1 U2573 ( .A(n12713), .B(n12959), .C(n1366), .Y(n5664) );
  NAND2X1 U2574 ( .A(ram[1227]), .B(n12959), .Y(n1366) );
  OAI21X1 U2575 ( .A(n12707), .B(n12959), .C(n1367), .Y(n5665) );
  NAND2X1 U2576 ( .A(ram[1228]), .B(n12959), .Y(n1367) );
  OAI21X1 U2577 ( .A(n12701), .B(n12959), .C(n1368), .Y(n5666) );
  NAND2X1 U2578 ( .A(ram[1229]), .B(n12959), .Y(n1368) );
  OAI21X1 U2579 ( .A(n12692), .B(n12959), .C(n1369), .Y(n5667) );
  NAND2X1 U2580 ( .A(ram[1230]), .B(n12959), .Y(n1369) );
  OAI21X1 U2581 ( .A(n12686), .B(n12959), .C(n1370), .Y(n5668) );
  NAND2X1 U2582 ( .A(ram[1231]), .B(n12959), .Y(n1370) );
  OAI21X1 U2584 ( .A(n12777), .B(n12958), .C(n1372), .Y(n5669) );
  NAND2X1 U2585 ( .A(ram[1232]), .B(n12958), .Y(n1372) );
  OAI21X1 U2586 ( .A(n12771), .B(n12958), .C(n1373), .Y(n5670) );
  NAND2X1 U2587 ( .A(ram[1233]), .B(n12958), .Y(n1373) );
  OAI21X1 U2588 ( .A(n12766), .B(n12958), .C(n1374), .Y(n5671) );
  NAND2X1 U2589 ( .A(ram[1234]), .B(n12958), .Y(n1374) );
  OAI21X1 U2590 ( .A(n12760), .B(n12958), .C(n1375), .Y(n5672) );
  NAND2X1 U2591 ( .A(ram[1235]), .B(n12958), .Y(n1375) );
  OAI21X1 U2592 ( .A(n12754), .B(n12958), .C(n1376), .Y(n5673) );
  NAND2X1 U2593 ( .A(ram[1236]), .B(n12958), .Y(n1376) );
  OAI21X1 U2594 ( .A(n12748), .B(n12958), .C(n1377), .Y(n5674) );
  NAND2X1 U2595 ( .A(ram[1237]), .B(n12958), .Y(n1377) );
  OAI21X1 U2596 ( .A(n12742), .B(n12958), .C(n1378), .Y(n5675) );
  NAND2X1 U2597 ( .A(ram[1238]), .B(n12958), .Y(n1378) );
  OAI21X1 U2598 ( .A(n12736), .B(n12958), .C(n1379), .Y(n5676) );
  NAND2X1 U2599 ( .A(ram[1239]), .B(n12958), .Y(n1379) );
  OAI21X1 U2600 ( .A(n12730), .B(n12958), .C(n1380), .Y(n5677) );
  NAND2X1 U2601 ( .A(ram[1240]), .B(n12958), .Y(n1380) );
  OAI21X1 U2602 ( .A(n12724), .B(n12958), .C(n1381), .Y(n5678) );
  NAND2X1 U2603 ( .A(ram[1241]), .B(n12958), .Y(n1381) );
  OAI21X1 U2604 ( .A(n12718), .B(n12958), .C(n1382), .Y(n5679) );
  NAND2X1 U2605 ( .A(ram[1242]), .B(n12958), .Y(n1382) );
  OAI21X1 U2606 ( .A(n12712), .B(n12958), .C(n1383), .Y(n5680) );
  NAND2X1 U2607 ( .A(ram[1243]), .B(n12958), .Y(n1383) );
  OAI21X1 U2608 ( .A(n12706), .B(n12958), .C(n1384), .Y(n5681) );
  NAND2X1 U2609 ( .A(ram[1244]), .B(n12958), .Y(n1384) );
  OAI21X1 U2610 ( .A(n12700), .B(n12958), .C(n1385), .Y(n5682) );
  NAND2X1 U2611 ( .A(ram[1245]), .B(n12958), .Y(n1385) );
  OAI21X1 U2612 ( .A(n12693), .B(n12958), .C(n1386), .Y(n5683) );
  NAND2X1 U2613 ( .A(ram[1246]), .B(n12958), .Y(n1386) );
  OAI21X1 U2614 ( .A(n12687), .B(n12958), .C(n1387), .Y(n5684) );
  NAND2X1 U2615 ( .A(ram[1247]), .B(n12958), .Y(n1387) );
  OAI21X1 U2617 ( .A(n12776), .B(n12957), .C(n1389), .Y(n5685) );
  NAND2X1 U2618 ( .A(ram[1248]), .B(n12957), .Y(n1389) );
  OAI21X1 U2619 ( .A(n12770), .B(n12957), .C(n1390), .Y(n5686) );
  NAND2X1 U2620 ( .A(ram[1249]), .B(n12957), .Y(n1390) );
  OAI21X1 U2621 ( .A(n12764), .B(n12957), .C(n1391), .Y(n5687) );
  NAND2X1 U2622 ( .A(ram[1250]), .B(n12957), .Y(n1391) );
  OAI21X1 U2623 ( .A(n12758), .B(n12957), .C(n1392), .Y(n5688) );
  NAND2X1 U2624 ( .A(ram[1251]), .B(n12957), .Y(n1392) );
  OAI21X1 U2625 ( .A(n12752), .B(n12957), .C(n1393), .Y(n5689) );
  NAND2X1 U2626 ( .A(ram[1252]), .B(n12957), .Y(n1393) );
  OAI21X1 U2627 ( .A(n12746), .B(n12957), .C(n1394), .Y(n5690) );
  NAND2X1 U2628 ( .A(ram[1253]), .B(n12957), .Y(n1394) );
  OAI21X1 U2629 ( .A(n12740), .B(n12957), .C(n1395), .Y(n5691) );
  NAND2X1 U2630 ( .A(ram[1254]), .B(n12957), .Y(n1395) );
  OAI21X1 U2631 ( .A(n12734), .B(n12957), .C(n1396), .Y(n5692) );
  NAND2X1 U2632 ( .A(ram[1255]), .B(n12957), .Y(n1396) );
  OAI21X1 U2633 ( .A(n12728), .B(n12957), .C(n1397), .Y(n5693) );
  NAND2X1 U2634 ( .A(ram[1256]), .B(n12957), .Y(n1397) );
  OAI21X1 U2635 ( .A(n12722), .B(n12957), .C(n1398), .Y(n5694) );
  NAND2X1 U2636 ( .A(ram[1257]), .B(n12957), .Y(n1398) );
  OAI21X1 U2637 ( .A(n12716), .B(n12957), .C(n1399), .Y(n5695) );
  NAND2X1 U2638 ( .A(ram[1258]), .B(n12957), .Y(n1399) );
  OAI21X1 U2639 ( .A(n12710), .B(n12957), .C(n1400), .Y(n5696) );
  NAND2X1 U2640 ( .A(ram[1259]), .B(n12957), .Y(n1400) );
  OAI21X1 U2641 ( .A(n12704), .B(n12957), .C(n1401), .Y(n5697) );
  NAND2X1 U2642 ( .A(ram[1260]), .B(n12957), .Y(n1401) );
  OAI21X1 U2643 ( .A(n12698), .B(n12957), .C(n1402), .Y(n5698) );
  NAND2X1 U2644 ( .A(ram[1261]), .B(n12957), .Y(n1402) );
  OAI21X1 U2645 ( .A(n12692), .B(n12957), .C(n1403), .Y(n5699) );
  NAND2X1 U2646 ( .A(ram[1262]), .B(n12957), .Y(n1403) );
  OAI21X1 U2647 ( .A(n12686), .B(n12957), .C(n1404), .Y(n5700) );
  NAND2X1 U2648 ( .A(ram[1263]), .B(n12957), .Y(n1404) );
  OAI21X1 U2650 ( .A(n12779), .B(n12956), .C(n1406), .Y(n5701) );
  NAND2X1 U2651 ( .A(ram[1264]), .B(n12956), .Y(n1406) );
  OAI21X1 U2652 ( .A(n12773), .B(n12956), .C(n1407), .Y(n5702) );
  NAND2X1 U2653 ( .A(ram[1265]), .B(n12956), .Y(n1407) );
  OAI21X1 U2654 ( .A(n12767), .B(n12956), .C(n1408), .Y(n5703) );
  NAND2X1 U2655 ( .A(ram[1266]), .B(n12956), .Y(n1408) );
  OAI21X1 U2656 ( .A(n12761), .B(n12956), .C(n1409), .Y(n5704) );
  NAND2X1 U2657 ( .A(ram[1267]), .B(n12956), .Y(n1409) );
  OAI21X1 U2658 ( .A(n12755), .B(n12956), .C(n1410), .Y(n5705) );
  NAND2X1 U2659 ( .A(ram[1268]), .B(n12956), .Y(n1410) );
  OAI21X1 U2660 ( .A(n12749), .B(n12956), .C(n1411), .Y(n5706) );
  NAND2X1 U2661 ( .A(ram[1269]), .B(n12956), .Y(n1411) );
  OAI21X1 U2662 ( .A(n12743), .B(n12956), .C(n1412), .Y(n5707) );
  NAND2X1 U2663 ( .A(ram[1270]), .B(n12956), .Y(n1412) );
  OAI21X1 U2664 ( .A(n12737), .B(n12956), .C(n1413), .Y(n5708) );
  NAND2X1 U2665 ( .A(ram[1271]), .B(n12956), .Y(n1413) );
  OAI21X1 U2666 ( .A(n12731), .B(n12956), .C(n1414), .Y(n5709) );
  NAND2X1 U2667 ( .A(ram[1272]), .B(n12956), .Y(n1414) );
  OAI21X1 U2668 ( .A(n12725), .B(n12956), .C(n1415), .Y(n5710) );
  NAND2X1 U2669 ( .A(ram[1273]), .B(n12956), .Y(n1415) );
  OAI21X1 U2670 ( .A(n12719), .B(n12956), .C(n1416), .Y(n5711) );
  NAND2X1 U2671 ( .A(ram[1274]), .B(n12956), .Y(n1416) );
  OAI21X1 U2672 ( .A(n12713), .B(n12956), .C(n1417), .Y(n5712) );
  NAND2X1 U2673 ( .A(ram[1275]), .B(n12956), .Y(n1417) );
  OAI21X1 U2674 ( .A(n12707), .B(n12956), .C(n1418), .Y(n5713) );
  NAND2X1 U2675 ( .A(ram[1276]), .B(n12956), .Y(n1418) );
  OAI21X1 U2676 ( .A(n12701), .B(n12956), .C(n1419), .Y(n5714) );
  NAND2X1 U2677 ( .A(ram[1277]), .B(n12956), .Y(n1419) );
  OAI21X1 U2678 ( .A(n12695), .B(n12956), .C(n1420), .Y(n5715) );
  NAND2X1 U2679 ( .A(ram[1278]), .B(n12956), .Y(n1420) );
  OAI21X1 U2680 ( .A(n12689), .B(n12956), .C(n1421), .Y(n5716) );
  NAND2X1 U2681 ( .A(ram[1279]), .B(n12956), .Y(n1421) );
  NAND3X1 U2683 ( .A(mem_write_en), .B(n327), .C(n1423), .Y(n1422) );
  OAI21X1 U2684 ( .A(n12778), .B(n12955), .C(n1425), .Y(n5717) );
  NAND2X1 U2685 ( .A(ram[1280]), .B(n12955), .Y(n1425) );
  OAI21X1 U2686 ( .A(n12772), .B(n12955), .C(n1426), .Y(n5718) );
  NAND2X1 U2687 ( .A(ram[1281]), .B(n12955), .Y(n1426) );
  OAI21X1 U2688 ( .A(n12766), .B(n12955), .C(n1427), .Y(n5719) );
  NAND2X1 U2689 ( .A(ram[1282]), .B(n12955), .Y(n1427) );
  OAI21X1 U2690 ( .A(n12760), .B(n12955), .C(n1428), .Y(n5720) );
  NAND2X1 U2691 ( .A(ram[1283]), .B(n12955), .Y(n1428) );
  OAI21X1 U2692 ( .A(n12754), .B(n12955), .C(n1429), .Y(n5721) );
  NAND2X1 U2693 ( .A(ram[1284]), .B(n12955), .Y(n1429) );
  OAI21X1 U2694 ( .A(n12748), .B(n12955), .C(n1430), .Y(n5722) );
  NAND2X1 U2695 ( .A(ram[1285]), .B(n12955), .Y(n1430) );
  OAI21X1 U2696 ( .A(n12742), .B(n12955), .C(n1431), .Y(n5723) );
  NAND2X1 U2697 ( .A(ram[1286]), .B(n12955), .Y(n1431) );
  OAI21X1 U2698 ( .A(n12736), .B(n12955), .C(n1432), .Y(n5724) );
  NAND2X1 U2699 ( .A(ram[1287]), .B(n12955), .Y(n1432) );
  OAI21X1 U2700 ( .A(n12730), .B(n12955), .C(n1433), .Y(n5725) );
  NAND2X1 U2701 ( .A(ram[1288]), .B(n12955), .Y(n1433) );
  OAI21X1 U2702 ( .A(n12724), .B(n12955), .C(n1434), .Y(n5726) );
  NAND2X1 U2703 ( .A(ram[1289]), .B(n12955), .Y(n1434) );
  OAI21X1 U2704 ( .A(n12718), .B(n12955), .C(n1435), .Y(n5727) );
  NAND2X1 U2705 ( .A(ram[1290]), .B(n12955), .Y(n1435) );
  OAI21X1 U2706 ( .A(n12712), .B(n12955), .C(n1436), .Y(n5728) );
  NAND2X1 U2707 ( .A(ram[1291]), .B(n12955), .Y(n1436) );
  OAI21X1 U2708 ( .A(n12706), .B(n12955), .C(n1437), .Y(n5729) );
  NAND2X1 U2709 ( .A(ram[1292]), .B(n12955), .Y(n1437) );
  OAI21X1 U2710 ( .A(n12700), .B(n12955), .C(n1438), .Y(n5730) );
  NAND2X1 U2711 ( .A(ram[1293]), .B(n12955), .Y(n1438) );
  OAI21X1 U2712 ( .A(n12694), .B(n12955), .C(n1439), .Y(n5731) );
  NAND2X1 U2713 ( .A(ram[1294]), .B(n12955), .Y(n1439) );
  OAI21X1 U2714 ( .A(n12688), .B(n12955), .C(n1440), .Y(n5732) );
  NAND2X1 U2715 ( .A(ram[1295]), .B(n12955), .Y(n1440) );
  OAI21X1 U2717 ( .A(n12777), .B(n12954), .C(n1442), .Y(n5733) );
  NAND2X1 U2718 ( .A(ram[1296]), .B(n12954), .Y(n1442) );
  OAI21X1 U2719 ( .A(n12771), .B(n12954), .C(n1443), .Y(n5734) );
  NAND2X1 U2720 ( .A(ram[1297]), .B(n12954), .Y(n1443) );
  OAI21X1 U2721 ( .A(n12765), .B(n12954), .C(n1444), .Y(n5735) );
  NAND2X1 U2722 ( .A(ram[1298]), .B(n12954), .Y(n1444) );
  OAI21X1 U2723 ( .A(n12759), .B(n12954), .C(n1445), .Y(n5736) );
  NAND2X1 U2724 ( .A(ram[1299]), .B(n12954), .Y(n1445) );
  OAI21X1 U2725 ( .A(n12753), .B(n12954), .C(n1446), .Y(n5737) );
  NAND2X1 U2726 ( .A(ram[1300]), .B(n12954), .Y(n1446) );
  OAI21X1 U2727 ( .A(n12747), .B(n12954), .C(n1447), .Y(n5738) );
  NAND2X1 U2728 ( .A(ram[1301]), .B(n12954), .Y(n1447) );
  OAI21X1 U2729 ( .A(n12741), .B(n12954), .C(n1448), .Y(n5739) );
  NAND2X1 U2730 ( .A(ram[1302]), .B(n12954), .Y(n1448) );
  OAI21X1 U2731 ( .A(n12735), .B(n12954), .C(n1449), .Y(n5740) );
  NAND2X1 U2732 ( .A(ram[1303]), .B(n12954), .Y(n1449) );
  OAI21X1 U2733 ( .A(n12729), .B(n12954), .C(n1450), .Y(n5741) );
  NAND2X1 U2734 ( .A(ram[1304]), .B(n12954), .Y(n1450) );
  OAI21X1 U2735 ( .A(n12723), .B(n12954), .C(n1451), .Y(n5742) );
  NAND2X1 U2736 ( .A(ram[1305]), .B(n12954), .Y(n1451) );
  OAI21X1 U2737 ( .A(n12717), .B(n12954), .C(n1452), .Y(n5743) );
  NAND2X1 U2738 ( .A(ram[1306]), .B(n12954), .Y(n1452) );
  OAI21X1 U2739 ( .A(n12711), .B(n12954), .C(n1453), .Y(n5744) );
  NAND2X1 U2740 ( .A(ram[1307]), .B(n12954), .Y(n1453) );
  OAI21X1 U2741 ( .A(n12705), .B(n12954), .C(n1454), .Y(n5745) );
  NAND2X1 U2742 ( .A(ram[1308]), .B(n12954), .Y(n1454) );
  OAI21X1 U2743 ( .A(n12699), .B(n12954), .C(n1455), .Y(n5746) );
  NAND2X1 U2744 ( .A(ram[1309]), .B(n12954), .Y(n1455) );
  OAI21X1 U2745 ( .A(n12693), .B(n12954), .C(n1456), .Y(n5747) );
  NAND2X1 U2746 ( .A(ram[1310]), .B(n12954), .Y(n1456) );
  OAI21X1 U2747 ( .A(n12687), .B(n12954), .C(n1457), .Y(n5748) );
  NAND2X1 U2748 ( .A(ram[1311]), .B(n12954), .Y(n1457) );
  OAI21X1 U2750 ( .A(n12775), .B(n12953), .C(n1459), .Y(n5749) );
  NAND2X1 U2751 ( .A(ram[1312]), .B(n12953), .Y(n1459) );
  OAI21X1 U2752 ( .A(n12769), .B(n12953), .C(n1460), .Y(n5750) );
  NAND2X1 U2753 ( .A(ram[1313]), .B(n12953), .Y(n1460) );
  OAI21X1 U2754 ( .A(n12767), .B(n12953), .C(n1461), .Y(n5751) );
  NAND2X1 U2755 ( .A(ram[1314]), .B(n12953), .Y(n1461) );
  OAI21X1 U2756 ( .A(n12761), .B(n12953), .C(n1462), .Y(n5752) );
  NAND2X1 U2757 ( .A(ram[1315]), .B(n12953), .Y(n1462) );
  OAI21X1 U2758 ( .A(n12755), .B(n12953), .C(n1463), .Y(n5753) );
  NAND2X1 U2759 ( .A(ram[1316]), .B(n12953), .Y(n1463) );
  OAI21X1 U2760 ( .A(n12749), .B(n12953), .C(n1464), .Y(n5754) );
  NAND2X1 U2761 ( .A(ram[1317]), .B(n12953), .Y(n1464) );
  OAI21X1 U2762 ( .A(n12743), .B(n12953), .C(n1465), .Y(n5755) );
  NAND2X1 U2763 ( .A(ram[1318]), .B(n12953), .Y(n1465) );
  OAI21X1 U2764 ( .A(n12737), .B(n12953), .C(n1466), .Y(n5756) );
  NAND2X1 U2765 ( .A(ram[1319]), .B(n12953), .Y(n1466) );
  OAI21X1 U2766 ( .A(n12731), .B(n12953), .C(n1467), .Y(n5757) );
  NAND2X1 U2767 ( .A(ram[1320]), .B(n12953), .Y(n1467) );
  OAI21X1 U2768 ( .A(n12725), .B(n12953), .C(n1468), .Y(n5758) );
  NAND2X1 U2769 ( .A(ram[1321]), .B(n12953), .Y(n1468) );
  OAI21X1 U2770 ( .A(n12719), .B(n12953), .C(n1469), .Y(n5759) );
  NAND2X1 U2771 ( .A(ram[1322]), .B(n12953), .Y(n1469) );
  OAI21X1 U2772 ( .A(n12713), .B(n12953), .C(n1470), .Y(n5760) );
  NAND2X1 U2773 ( .A(ram[1323]), .B(n12953), .Y(n1470) );
  OAI21X1 U2774 ( .A(n12707), .B(n12953), .C(n1471), .Y(n5761) );
  NAND2X1 U2775 ( .A(ram[1324]), .B(n12953), .Y(n1471) );
  OAI21X1 U2776 ( .A(n12701), .B(n12953), .C(n1472), .Y(n5762) );
  NAND2X1 U2777 ( .A(ram[1325]), .B(n12953), .Y(n1472) );
  OAI21X1 U2778 ( .A(n12691), .B(n12953), .C(n1473), .Y(n5763) );
  NAND2X1 U2779 ( .A(ram[1326]), .B(n12953), .Y(n1473) );
  OAI21X1 U2780 ( .A(n12685), .B(n12953), .C(n1474), .Y(n5764) );
  NAND2X1 U2781 ( .A(ram[1327]), .B(n12953), .Y(n1474) );
  OAI21X1 U2783 ( .A(n12775), .B(n12952), .C(n1476), .Y(n5765) );
  NAND2X1 U2784 ( .A(ram[1328]), .B(n12952), .Y(n1476) );
  OAI21X1 U2785 ( .A(n12769), .B(n12952), .C(n1477), .Y(n5766) );
  NAND2X1 U2786 ( .A(ram[1329]), .B(n12952), .Y(n1477) );
  OAI21X1 U2787 ( .A(n12766), .B(n12952), .C(n1478), .Y(n5767) );
  NAND2X1 U2788 ( .A(ram[1330]), .B(n12952), .Y(n1478) );
  OAI21X1 U2789 ( .A(n12760), .B(n12952), .C(n1479), .Y(n5768) );
  NAND2X1 U2790 ( .A(ram[1331]), .B(n12952), .Y(n1479) );
  OAI21X1 U2791 ( .A(n12754), .B(n12952), .C(n1480), .Y(n5769) );
  NAND2X1 U2792 ( .A(ram[1332]), .B(n12952), .Y(n1480) );
  OAI21X1 U2793 ( .A(n12748), .B(n12952), .C(n1481), .Y(n5770) );
  NAND2X1 U2794 ( .A(ram[1333]), .B(n12952), .Y(n1481) );
  OAI21X1 U2795 ( .A(n12742), .B(n12952), .C(n1482), .Y(n5771) );
  NAND2X1 U2796 ( .A(ram[1334]), .B(n12952), .Y(n1482) );
  OAI21X1 U2797 ( .A(n12736), .B(n12952), .C(n1483), .Y(n5772) );
  NAND2X1 U2798 ( .A(ram[1335]), .B(n12952), .Y(n1483) );
  OAI21X1 U2799 ( .A(n12730), .B(n12952), .C(n1484), .Y(n5773) );
  NAND2X1 U2800 ( .A(ram[1336]), .B(n12952), .Y(n1484) );
  OAI21X1 U2801 ( .A(n12724), .B(n12952), .C(n1485), .Y(n5774) );
  NAND2X1 U2802 ( .A(ram[1337]), .B(n12952), .Y(n1485) );
  OAI21X1 U2803 ( .A(n12718), .B(n12952), .C(n1486), .Y(n5775) );
  NAND2X1 U2804 ( .A(ram[1338]), .B(n12952), .Y(n1486) );
  OAI21X1 U2805 ( .A(n12712), .B(n12952), .C(n1487), .Y(n5776) );
  NAND2X1 U2806 ( .A(ram[1339]), .B(n12952), .Y(n1487) );
  OAI21X1 U2807 ( .A(n12706), .B(n12952), .C(n1488), .Y(n5777) );
  NAND2X1 U2808 ( .A(ram[1340]), .B(n12952), .Y(n1488) );
  OAI21X1 U2809 ( .A(n12700), .B(n12952), .C(n1489), .Y(n5778) );
  NAND2X1 U2810 ( .A(ram[1341]), .B(n12952), .Y(n1489) );
  OAI21X1 U2811 ( .A(n12691), .B(n12952), .C(n1490), .Y(n5779) );
  NAND2X1 U2812 ( .A(ram[1342]), .B(n12952), .Y(n1490) );
  OAI21X1 U2813 ( .A(n12685), .B(n12952), .C(n1491), .Y(n5780) );
  NAND2X1 U2814 ( .A(ram[1343]), .B(n12952), .Y(n1491) );
  OAI21X1 U2816 ( .A(n12779), .B(n12951), .C(n1493), .Y(n5781) );
  NAND2X1 U2817 ( .A(ram[1344]), .B(n12951), .Y(n1493) );
  OAI21X1 U2818 ( .A(n12773), .B(n12951), .C(n1494), .Y(n5782) );
  NAND2X1 U2819 ( .A(ram[1345]), .B(n12951), .Y(n1494) );
  OAI21X1 U2820 ( .A(n12765), .B(n12951), .C(n1495), .Y(n5783) );
  NAND2X1 U2821 ( .A(ram[1346]), .B(n12951), .Y(n1495) );
  OAI21X1 U2822 ( .A(n12759), .B(n12951), .C(n1496), .Y(n5784) );
  NAND2X1 U2823 ( .A(ram[1347]), .B(n12951), .Y(n1496) );
  OAI21X1 U2824 ( .A(n12753), .B(n12951), .C(n1497), .Y(n5785) );
  NAND2X1 U2825 ( .A(ram[1348]), .B(n12951), .Y(n1497) );
  OAI21X1 U2826 ( .A(n12747), .B(n12951), .C(n1498), .Y(n5786) );
  NAND2X1 U2827 ( .A(ram[1349]), .B(n12951), .Y(n1498) );
  OAI21X1 U2828 ( .A(n12741), .B(n12951), .C(n1499), .Y(n5787) );
  NAND2X1 U2829 ( .A(ram[1350]), .B(n12951), .Y(n1499) );
  OAI21X1 U2830 ( .A(n12735), .B(n12951), .C(n1500), .Y(n5788) );
  NAND2X1 U2831 ( .A(ram[1351]), .B(n12951), .Y(n1500) );
  OAI21X1 U2832 ( .A(n12729), .B(n12951), .C(n1501), .Y(n5789) );
  NAND2X1 U2833 ( .A(ram[1352]), .B(n12951), .Y(n1501) );
  OAI21X1 U2834 ( .A(n12723), .B(n12951), .C(n1502), .Y(n5790) );
  NAND2X1 U2835 ( .A(ram[1353]), .B(n12951), .Y(n1502) );
  OAI21X1 U2836 ( .A(n12717), .B(n12951), .C(n1503), .Y(n5791) );
  NAND2X1 U2837 ( .A(ram[1354]), .B(n12951), .Y(n1503) );
  OAI21X1 U2838 ( .A(n12711), .B(n12951), .C(n1504), .Y(n5792) );
  NAND2X1 U2839 ( .A(ram[1355]), .B(n12951), .Y(n1504) );
  OAI21X1 U2840 ( .A(n12705), .B(n12951), .C(n1505), .Y(n5793) );
  NAND2X1 U2841 ( .A(ram[1356]), .B(n12951), .Y(n1505) );
  OAI21X1 U2842 ( .A(n12699), .B(n12951), .C(n1506), .Y(n5794) );
  NAND2X1 U2843 ( .A(ram[1357]), .B(n12951), .Y(n1506) );
  OAI21X1 U2844 ( .A(n12695), .B(n12951), .C(n1507), .Y(n5795) );
  NAND2X1 U2845 ( .A(ram[1358]), .B(n12951), .Y(n1507) );
  OAI21X1 U2846 ( .A(n12689), .B(n12951), .C(n1508), .Y(n5796) );
  NAND2X1 U2847 ( .A(ram[1359]), .B(n12951), .Y(n1508) );
  OAI21X1 U2849 ( .A(n12778), .B(n12950), .C(n1510), .Y(n5797) );
  NAND2X1 U2850 ( .A(ram[1360]), .B(n12950), .Y(n1510) );
  OAI21X1 U2851 ( .A(n12772), .B(n12950), .C(n1511), .Y(n5798) );
  NAND2X1 U2852 ( .A(ram[1361]), .B(n12950), .Y(n1511) );
  OAI21X1 U2853 ( .A(n12763), .B(n12950), .C(n1512), .Y(n5799) );
  NAND2X1 U2854 ( .A(ram[1362]), .B(n12950), .Y(n1512) );
  OAI21X1 U2855 ( .A(n12757), .B(n12950), .C(n1513), .Y(n5800) );
  NAND2X1 U2856 ( .A(ram[1363]), .B(n12950), .Y(n1513) );
  OAI21X1 U2857 ( .A(n12751), .B(n12950), .C(n1514), .Y(n5801) );
  NAND2X1 U2858 ( .A(ram[1364]), .B(n12950), .Y(n1514) );
  OAI21X1 U2859 ( .A(n12745), .B(n12950), .C(n1515), .Y(n5802) );
  NAND2X1 U2860 ( .A(ram[1365]), .B(n12950), .Y(n1515) );
  OAI21X1 U2861 ( .A(n12739), .B(n12950), .C(n1516), .Y(n5803) );
  NAND2X1 U2862 ( .A(ram[1366]), .B(n12950), .Y(n1516) );
  OAI21X1 U2863 ( .A(n12733), .B(n12950), .C(n1517), .Y(n5804) );
  NAND2X1 U2864 ( .A(ram[1367]), .B(n12950), .Y(n1517) );
  OAI21X1 U2865 ( .A(n12727), .B(n12950), .C(n1518), .Y(n5805) );
  NAND2X1 U2866 ( .A(ram[1368]), .B(n12950), .Y(n1518) );
  OAI21X1 U2867 ( .A(n12721), .B(n12950), .C(n1519), .Y(n5806) );
  NAND2X1 U2868 ( .A(ram[1369]), .B(n12950), .Y(n1519) );
  OAI21X1 U2869 ( .A(n12715), .B(n12950), .C(n1520), .Y(n5807) );
  NAND2X1 U2870 ( .A(ram[1370]), .B(n12950), .Y(n1520) );
  OAI21X1 U2871 ( .A(n12709), .B(n12950), .C(n1521), .Y(n5808) );
  NAND2X1 U2872 ( .A(ram[1371]), .B(n12950), .Y(n1521) );
  OAI21X1 U2873 ( .A(n12703), .B(n12950), .C(n1522), .Y(n5809) );
  NAND2X1 U2874 ( .A(ram[1372]), .B(n12950), .Y(n1522) );
  OAI21X1 U2875 ( .A(n12697), .B(n12950), .C(n1523), .Y(n5810) );
  NAND2X1 U2876 ( .A(ram[1373]), .B(n12950), .Y(n1523) );
  OAI21X1 U2877 ( .A(n12694), .B(n12950), .C(n1524), .Y(n5811) );
  NAND2X1 U2878 ( .A(ram[1374]), .B(n12950), .Y(n1524) );
  OAI21X1 U2879 ( .A(n12688), .B(n12950), .C(n1525), .Y(n5812) );
  NAND2X1 U2880 ( .A(ram[1375]), .B(n12950), .Y(n1525) );
  OAI21X1 U2882 ( .A(n12777), .B(n12949), .C(n1527), .Y(n5813) );
  NAND2X1 U2883 ( .A(ram[1376]), .B(n12949), .Y(n1527) );
  OAI21X1 U2884 ( .A(n12771), .B(n12949), .C(n1528), .Y(n5814) );
  NAND2X1 U2885 ( .A(ram[1377]), .B(n12949), .Y(n1528) );
  OAI21X1 U2886 ( .A(n12764), .B(n12949), .C(n1529), .Y(n5815) );
  NAND2X1 U2887 ( .A(ram[1378]), .B(n12949), .Y(n1529) );
  OAI21X1 U2888 ( .A(n12758), .B(n12949), .C(n1530), .Y(n5816) );
  NAND2X1 U2889 ( .A(ram[1379]), .B(n12949), .Y(n1530) );
  OAI21X1 U2890 ( .A(n12752), .B(n12949), .C(n1531), .Y(n5817) );
  NAND2X1 U2891 ( .A(ram[1380]), .B(n12949), .Y(n1531) );
  OAI21X1 U2892 ( .A(n12746), .B(n12949), .C(n1532), .Y(n5818) );
  NAND2X1 U2893 ( .A(ram[1381]), .B(n12949), .Y(n1532) );
  OAI21X1 U2894 ( .A(n12740), .B(n12949), .C(n1533), .Y(n5819) );
  NAND2X1 U2895 ( .A(ram[1382]), .B(n12949), .Y(n1533) );
  OAI21X1 U2896 ( .A(n12734), .B(n12949), .C(n1534), .Y(n5820) );
  NAND2X1 U2897 ( .A(ram[1383]), .B(n12949), .Y(n1534) );
  OAI21X1 U2898 ( .A(n12728), .B(n12949), .C(n1535), .Y(n5821) );
  NAND2X1 U2899 ( .A(ram[1384]), .B(n12949), .Y(n1535) );
  OAI21X1 U2900 ( .A(n12722), .B(n12949), .C(n1536), .Y(n5822) );
  NAND2X1 U2901 ( .A(ram[1385]), .B(n12949), .Y(n1536) );
  OAI21X1 U2902 ( .A(n12716), .B(n12949), .C(n1537), .Y(n5823) );
  NAND2X1 U2903 ( .A(ram[1386]), .B(n12949), .Y(n1537) );
  OAI21X1 U2904 ( .A(n12710), .B(n12949), .C(n1538), .Y(n5824) );
  NAND2X1 U2905 ( .A(ram[1387]), .B(n12949), .Y(n1538) );
  OAI21X1 U2906 ( .A(n12704), .B(n12949), .C(n1539), .Y(n5825) );
  NAND2X1 U2907 ( .A(ram[1388]), .B(n12949), .Y(n1539) );
  OAI21X1 U2908 ( .A(n12698), .B(n12949), .C(n1540), .Y(n5826) );
  NAND2X1 U2909 ( .A(ram[1389]), .B(n12949), .Y(n1540) );
  OAI21X1 U2910 ( .A(n12693), .B(n12949), .C(n1541), .Y(n5827) );
  NAND2X1 U2911 ( .A(ram[1390]), .B(n12949), .Y(n1541) );
  OAI21X1 U2912 ( .A(n12687), .B(n12949), .C(n1542), .Y(n5828) );
  NAND2X1 U2913 ( .A(ram[1391]), .B(n12949), .Y(n1542) );
  OAI21X1 U2915 ( .A(n12776), .B(n12948), .C(n1544), .Y(n5829) );
  NAND2X1 U2916 ( .A(ram[1392]), .B(n12948), .Y(n1544) );
  OAI21X1 U2917 ( .A(n12770), .B(n12948), .C(n1545), .Y(n5830) );
  NAND2X1 U2918 ( .A(ram[1393]), .B(n12948), .Y(n1545) );
  OAI21X1 U2919 ( .A(n12764), .B(n12948), .C(n1546), .Y(n5831) );
  NAND2X1 U2920 ( .A(ram[1394]), .B(n12948), .Y(n1546) );
  OAI21X1 U2921 ( .A(n12758), .B(n12948), .C(n1547), .Y(n5832) );
  NAND2X1 U2922 ( .A(ram[1395]), .B(n12948), .Y(n1547) );
  OAI21X1 U2923 ( .A(n12752), .B(n12948), .C(n1548), .Y(n5833) );
  NAND2X1 U2924 ( .A(ram[1396]), .B(n12948), .Y(n1548) );
  OAI21X1 U2925 ( .A(n12746), .B(n12948), .C(n1549), .Y(n5834) );
  NAND2X1 U2926 ( .A(ram[1397]), .B(n12948), .Y(n1549) );
  OAI21X1 U2927 ( .A(n12740), .B(n12948), .C(n1550), .Y(n5835) );
  NAND2X1 U2928 ( .A(ram[1398]), .B(n12948), .Y(n1550) );
  OAI21X1 U2929 ( .A(n12734), .B(n12948), .C(n1551), .Y(n5836) );
  NAND2X1 U2930 ( .A(ram[1399]), .B(n12948), .Y(n1551) );
  OAI21X1 U2931 ( .A(n12728), .B(n12948), .C(n1552), .Y(n5837) );
  NAND2X1 U2932 ( .A(ram[1400]), .B(n12948), .Y(n1552) );
  OAI21X1 U2933 ( .A(n12722), .B(n12948), .C(n1553), .Y(n5838) );
  NAND2X1 U2934 ( .A(ram[1401]), .B(n12948), .Y(n1553) );
  OAI21X1 U2935 ( .A(n12716), .B(n12948), .C(n1554), .Y(n5839) );
  NAND2X1 U2936 ( .A(ram[1402]), .B(n12948), .Y(n1554) );
  OAI21X1 U2937 ( .A(n12710), .B(n12948), .C(n1555), .Y(n5840) );
  NAND2X1 U2938 ( .A(ram[1403]), .B(n12948), .Y(n1555) );
  OAI21X1 U2939 ( .A(n12704), .B(n12948), .C(n1556), .Y(n5841) );
  NAND2X1 U2940 ( .A(ram[1404]), .B(n12948), .Y(n1556) );
  OAI21X1 U2941 ( .A(n12698), .B(n12948), .C(n1557), .Y(n5842) );
  NAND2X1 U2942 ( .A(ram[1405]), .B(n12948), .Y(n1557) );
  OAI21X1 U2943 ( .A(n12692), .B(n12948), .C(n1558), .Y(n5843) );
  NAND2X1 U2944 ( .A(ram[1406]), .B(n12948), .Y(n1558) );
  OAI21X1 U2945 ( .A(n12686), .B(n12948), .C(n1559), .Y(n5844) );
  NAND2X1 U2946 ( .A(ram[1407]), .B(n12948), .Y(n1559) );
  OAI21X1 U2948 ( .A(n12778), .B(n12947), .C(n1561), .Y(n5845) );
  NAND2X1 U2949 ( .A(ram[1408]), .B(n12947), .Y(n1561) );
  OAI21X1 U2950 ( .A(n12772), .B(n12947), .C(n1562), .Y(n5846) );
  NAND2X1 U2951 ( .A(ram[1409]), .B(n12947), .Y(n1562) );
  OAI21X1 U2952 ( .A(n12764), .B(n12947), .C(n1563), .Y(n5847) );
  NAND2X1 U2953 ( .A(ram[1410]), .B(n12947), .Y(n1563) );
  OAI21X1 U2954 ( .A(n12758), .B(n12947), .C(n1564), .Y(n5848) );
  NAND2X1 U2955 ( .A(ram[1411]), .B(n12947), .Y(n1564) );
  OAI21X1 U2956 ( .A(n12752), .B(n12947), .C(n1565), .Y(n5849) );
  NAND2X1 U2957 ( .A(ram[1412]), .B(n12947), .Y(n1565) );
  OAI21X1 U2958 ( .A(n12746), .B(n12947), .C(n1566), .Y(n5850) );
  NAND2X1 U2959 ( .A(ram[1413]), .B(n12947), .Y(n1566) );
  OAI21X1 U2960 ( .A(n12740), .B(n12947), .C(n1567), .Y(n5851) );
  NAND2X1 U2961 ( .A(ram[1414]), .B(n12947), .Y(n1567) );
  OAI21X1 U2962 ( .A(n12734), .B(n12947), .C(n1568), .Y(n5852) );
  NAND2X1 U2963 ( .A(ram[1415]), .B(n12947), .Y(n1568) );
  OAI21X1 U2964 ( .A(n12728), .B(n12947), .C(n1569), .Y(n5853) );
  NAND2X1 U2965 ( .A(ram[1416]), .B(n12947), .Y(n1569) );
  OAI21X1 U2966 ( .A(n12722), .B(n12947), .C(n1570), .Y(n5854) );
  NAND2X1 U2967 ( .A(ram[1417]), .B(n12947), .Y(n1570) );
  OAI21X1 U2968 ( .A(n12716), .B(n12947), .C(n1571), .Y(n5855) );
  NAND2X1 U2969 ( .A(ram[1418]), .B(n12947), .Y(n1571) );
  OAI21X1 U2970 ( .A(n12710), .B(n12947), .C(n1572), .Y(n5856) );
  NAND2X1 U2971 ( .A(ram[1419]), .B(n12947), .Y(n1572) );
  OAI21X1 U2972 ( .A(n12704), .B(n12947), .C(n1573), .Y(n5857) );
  NAND2X1 U2973 ( .A(ram[1420]), .B(n12947), .Y(n1573) );
  OAI21X1 U2974 ( .A(n12698), .B(n12947), .C(n1574), .Y(n5858) );
  NAND2X1 U2975 ( .A(ram[1421]), .B(n12947), .Y(n1574) );
  OAI21X1 U2976 ( .A(n12694), .B(n12947), .C(n1575), .Y(n5859) );
  NAND2X1 U2977 ( .A(ram[1422]), .B(n12947), .Y(n1575) );
  OAI21X1 U2978 ( .A(n12688), .B(n12947), .C(n1576), .Y(n5860) );
  NAND2X1 U2979 ( .A(ram[1423]), .B(n12947), .Y(n1576) );
  OAI21X1 U2981 ( .A(n12777), .B(n12946), .C(n1578), .Y(n5861) );
  NAND2X1 U2982 ( .A(ram[1424]), .B(n12946), .Y(n1578) );
  OAI21X1 U2983 ( .A(n12771), .B(n12946), .C(n1579), .Y(n5862) );
  NAND2X1 U2984 ( .A(ram[1425]), .B(n12946), .Y(n1579) );
  OAI21X1 U2985 ( .A(n12767), .B(n12946), .C(n1580), .Y(n5863) );
  NAND2X1 U2986 ( .A(ram[1426]), .B(n12946), .Y(n1580) );
  OAI21X1 U2987 ( .A(n12761), .B(n12946), .C(n1581), .Y(n5864) );
  NAND2X1 U2988 ( .A(ram[1427]), .B(n12946), .Y(n1581) );
  OAI21X1 U2989 ( .A(n12755), .B(n12946), .C(n1582), .Y(n5865) );
  NAND2X1 U2990 ( .A(ram[1428]), .B(n12946), .Y(n1582) );
  OAI21X1 U2991 ( .A(n12749), .B(n12946), .C(n1583), .Y(n5866) );
  NAND2X1 U2992 ( .A(ram[1429]), .B(n12946), .Y(n1583) );
  OAI21X1 U2993 ( .A(n12743), .B(n12946), .C(n1584), .Y(n5867) );
  NAND2X1 U2994 ( .A(ram[1430]), .B(n12946), .Y(n1584) );
  OAI21X1 U2995 ( .A(n12737), .B(n12946), .C(n1585), .Y(n5868) );
  NAND2X1 U2996 ( .A(ram[1431]), .B(n12946), .Y(n1585) );
  OAI21X1 U2997 ( .A(n12731), .B(n12946), .C(n1586), .Y(n5869) );
  NAND2X1 U2998 ( .A(ram[1432]), .B(n12946), .Y(n1586) );
  OAI21X1 U2999 ( .A(n12725), .B(n12946), .C(n1587), .Y(n5870) );
  NAND2X1 U3000 ( .A(ram[1433]), .B(n12946), .Y(n1587) );
  OAI21X1 U3001 ( .A(n12719), .B(n12946), .C(n1588), .Y(n5871) );
  NAND2X1 U3002 ( .A(ram[1434]), .B(n12946), .Y(n1588) );
  OAI21X1 U3003 ( .A(n12713), .B(n12946), .C(n1589), .Y(n5872) );
  NAND2X1 U3004 ( .A(ram[1435]), .B(n12946), .Y(n1589) );
  OAI21X1 U3005 ( .A(n12707), .B(n12946), .C(n1590), .Y(n5873) );
  NAND2X1 U3006 ( .A(ram[1436]), .B(n12946), .Y(n1590) );
  OAI21X1 U3007 ( .A(n12701), .B(n12946), .C(n1591), .Y(n5874) );
  NAND2X1 U3008 ( .A(ram[1437]), .B(n12946), .Y(n1591) );
  OAI21X1 U3009 ( .A(n12693), .B(n12946), .C(n1592), .Y(n5875) );
  NAND2X1 U3010 ( .A(ram[1438]), .B(n12946), .Y(n1592) );
  OAI21X1 U3011 ( .A(n12687), .B(n12946), .C(n1593), .Y(n5876) );
  NAND2X1 U3012 ( .A(ram[1439]), .B(n12946), .Y(n1593) );
  OAI21X1 U3014 ( .A(n12776), .B(n12945), .C(n1595), .Y(n5877) );
  NAND2X1 U3015 ( .A(ram[1440]), .B(n12945), .Y(n1595) );
  OAI21X1 U3016 ( .A(n12770), .B(n12945), .C(n1596), .Y(n5878) );
  NAND2X1 U3017 ( .A(ram[1441]), .B(n12945), .Y(n1596) );
  OAI21X1 U3018 ( .A(n12763), .B(n12945), .C(n1597), .Y(n5879) );
  NAND2X1 U3019 ( .A(ram[1442]), .B(n12945), .Y(n1597) );
  OAI21X1 U3020 ( .A(n12757), .B(n12945), .C(n1598), .Y(n5880) );
  NAND2X1 U3021 ( .A(ram[1443]), .B(n12945), .Y(n1598) );
  OAI21X1 U3022 ( .A(n12751), .B(n12945), .C(n1599), .Y(n5881) );
  NAND2X1 U3023 ( .A(ram[1444]), .B(n12945), .Y(n1599) );
  OAI21X1 U3024 ( .A(n12745), .B(n12945), .C(n1600), .Y(n5882) );
  NAND2X1 U3025 ( .A(ram[1445]), .B(n12945), .Y(n1600) );
  OAI21X1 U3026 ( .A(n12739), .B(n12945), .C(n1601), .Y(n5883) );
  NAND2X1 U3027 ( .A(ram[1446]), .B(n12945), .Y(n1601) );
  OAI21X1 U3028 ( .A(n12733), .B(n12945), .C(n1602), .Y(n5884) );
  NAND2X1 U3029 ( .A(ram[1447]), .B(n12945), .Y(n1602) );
  OAI21X1 U3030 ( .A(n12727), .B(n12945), .C(n1603), .Y(n5885) );
  NAND2X1 U3031 ( .A(ram[1448]), .B(n12945), .Y(n1603) );
  OAI21X1 U3032 ( .A(n12721), .B(n12945), .C(n1604), .Y(n5886) );
  NAND2X1 U3033 ( .A(ram[1449]), .B(n12945), .Y(n1604) );
  OAI21X1 U3034 ( .A(n12715), .B(n12945), .C(n1605), .Y(n5887) );
  NAND2X1 U3035 ( .A(ram[1450]), .B(n12945), .Y(n1605) );
  OAI21X1 U3036 ( .A(n12709), .B(n12945), .C(n1606), .Y(n5888) );
  NAND2X1 U3037 ( .A(ram[1451]), .B(n12945), .Y(n1606) );
  OAI21X1 U3038 ( .A(n12703), .B(n12945), .C(n1607), .Y(n5889) );
  NAND2X1 U3039 ( .A(ram[1452]), .B(n12945), .Y(n1607) );
  OAI21X1 U3040 ( .A(n12697), .B(n12945), .C(n1608), .Y(n5890) );
  NAND2X1 U3041 ( .A(ram[1453]), .B(n12945), .Y(n1608) );
  OAI21X1 U3042 ( .A(n12692), .B(n12945), .C(n1609), .Y(n5891) );
  NAND2X1 U3043 ( .A(ram[1454]), .B(n12945), .Y(n1609) );
  OAI21X1 U3044 ( .A(n12686), .B(n12945), .C(n1610), .Y(n5892) );
  NAND2X1 U3045 ( .A(ram[1455]), .B(n12945), .Y(n1610) );
  OAI21X1 U3047 ( .A(n12774), .B(n12944), .C(n1612), .Y(n5893) );
  NAND2X1 U3048 ( .A(ram[1456]), .B(n12944), .Y(n1612) );
  OAI21X1 U3049 ( .A(n12768), .B(n12944), .C(n1613), .Y(n5894) );
  NAND2X1 U3050 ( .A(ram[1457]), .B(n12944), .Y(n1613) );
  OAI21X1 U3051 ( .A(n12763), .B(n12944), .C(n1614), .Y(n5895) );
  NAND2X1 U3052 ( .A(ram[1458]), .B(n12944), .Y(n1614) );
  OAI21X1 U3053 ( .A(n12757), .B(n12944), .C(n1615), .Y(n5896) );
  NAND2X1 U3054 ( .A(ram[1459]), .B(n12944), .Y(n1615) );
  OAI21X1 U3055 ( .A(n12751), .B(n12944), .C(n1616), .Y(n5897) );
  NAND2X1 U3056 ( .A(ram[1460]), .B(n12944), .Y(n1616) );
  OAI21X1 U3057 ( .A(n12745), .B(n12944), .C(n1617), .Y(n5898) );
  NAND2X1 U3058 ( .A(ram[1461]), .B(n12944), .Y(n1617) );
  OAI21X1 U3059 ( .A(n12739), .B(n12944), .C(n1618), .Y(n5899) );
  NAND2X1 U3060 ( .A(ram[1462]), .B(n12944), .Y(n1618) );
  OAI21X1 U3061 ( .A(n12733), .B(n12944), .C(n1619), .Y(n5900) );
  NAND2X1 U3062 ( .A(ram[1463]), .B(n12944), .Y(n1619) );
  OAI21X1 U3063 ( .A(n12727), .B(n12944), .C(n1620), .Y(n5901) );
  NAND2X1 U3064 ( .A(ram[1464]), .B(n12944), .Y(n1620) );
  OAI21X1 U3065 ( .A(n12721), .B(n12944), .C(n1621), .Y(n5902) );
  NAND2X1 U3066 ( .A(ram[1465]), .B(n12944), .Y(n1621) );
  OAI21X1 U3067 ( .A(n12715), .B(n12944), .C(n1622), .Y(n5903) );
  NAND2X1 U3068 ( .A(ram[1466]), .B(n12944), .Y(n1622) );
  OAI21X1 U3069 ( .A(n12709), .B(n12944), .C(n1623), .Y(n5904) );
  NAND2X1 U3070 ( .A(ram[1467]), .B(n12944), .Y(n1623) );
  OAI21X1 U3071 ( .A(n12703), .B(n12944), .C(n1624), .Y(n5905) );
  NAND2X1 U3072 ( .A(ram[1468]), .B(n12944), .Y(n1624) );
  OAI21X1 U3073 ( .A(n12697), .B(n12944), .C(n1625), .Y(n5906) );
  NAND2X1 U3074 ( .A(ram[1469]), .B(n12944), .Y(n1625) );
  OAI21X1 U3075 ( .A(n12690), .B(n12944), .C(n1626), .Y(n5907) );
  NAND2X1 U3076 ( .A(ram[1470]), .B(n12944), .Y(n1626) );
  OAI21X1 U3077 ( .A(n12684), .B(n12944), .C(n1627), .Y(n5908) );
  NAND2X1 U3078 ( .A(ram[1471]), .B(n12944), .Y(n1627) );
  OAI21X1 U3080 ( .A(n12775), .B(n12943), .C(n1629), .Y(n5909) );
  NAND2X1 U3081 ( .A(ram[1472]), .B(n12943), .Y(n1629) );
  OAI21X1 U3082 ( .A(n12769), .B(n12943), .C(n1630), .Y(n5910) );
  NAND2X1 U3083 ( .A(ram[1473]), .B(n12943), .Y(n1630) );
  OAI21X1 U3084 ( .A(n13069), .B(n12943), .C(n1631), .Y(n5911) );
  NAND2X1 U3085 ( .A(ram[1474]), .B(n12943), .Y(n1631) );
  OAI21X1 U3086 ( .A(n13068), .B(n12943), .C(n1632), .Y(n5912) );
  NAND2X1 U3087 ( .A(ram[1475]), .B(n12943), .Y(n1632) );
  OAI21X1 U3088 ( .A(n13067), .B(n12943), .C(n1633), .Y(n5913) );
  NAND2X1 U3089 ( .A(ram[1476]), .B(n12943), .Y(n1633) );
  OAI21X1 U3090 ( .A(n13066), .B(n12943), .C(n1634), .Y(n5914) );
  NAND2X1 U3091 ( .A(ram[1477]), .B(n12943), .Y(n1634) );
  OAI21X1 U3092 ( .A(n13065), .B(n12943), .C(n1635), .Y(n5915) );
  NAND2X1 U3093 ( .A(ram[1478]), .B(n12943), .Y(n1635) );
  OAI21X1 U3094 ( .A(n13064), .B(n12943), .C(n1636), .Y(n5916) );
  NAND2X1 U3095 ( .A(ram[1479]), .B(n12943), .Y(n1636) );
  OAI21X1 U3096 ( .A(n13063), .B(n12943), .C(n1637), .Y(n5917) );
  NAND2X1 U3097 ( .A(ram[1480]), .B(n12943), .Y(n1637) );
  OAI21X1 U3098 ( .A(n13062), .B(n12943), .C(n1638), .Y(n5918) );
  NAND2X1 U3099 ( .A(ram[1481]), .B(n12943), .Y(n1638) );
  OAI21X1 U3100 ( .A(n13061), .B(n12943), .C(n1639), .Y(n5919) );
  NAND2X1 U3101 ( .A(ram[1482]), .B(n12943), .Y(n1639) );
  OAI21X1 U3102 ( .A(n13060), .B(n12943), .C(n1640), .Y(n5920) );
  NAND2X1 U3103 ( .A(ram[1483]), .B(n12943), .Y(n1640) );
  OAI21X1 U3104 ( .A(n13059), .B(n12943), .C(n1641), .Y(n5921) );
  NAND2X1 U3105 ( .A(ram[1484]), .B(n12943), .Y(n1641) );
  OAI21X1 U3106 ( .A(n13058), .B(n12943), .C(n1642), .Y(n5922) );
  NAND2X1 U3107 ( .A(ram[1485]), .B(n12943), .Y(n1642) );
  OAI21X1 U3108 ( .A(n12691), .B(n12943), .C(n1643), .Y(n5923) );
  NAND2X1 U3109 ( .A(ram[1486]), .B(n12943), .Y(n1643) );
  OAI21X1 U3110 ( .A(n12685), .B(n12943), .C(n1644), .Y(n5924) );
  NAND2X1 U3111 ( .A(ram[1487]), .B(n12943), .Y(n1644) );
  OAI21X1 U3113 ( .A(n12779), .B(n12942), .C(n1646), .Y(n5925) );
  NAND2X1 U3114 ( .A(ram[1488]), .B(n12942), .Y(n1646) );
  OAI21X1 U3115 ( .A(n12773), .B(n12942), .C(n1647), .Y(n5926) );
  NAND2X1 U3116 ( .A(ram[1489]), .B(n12942), .Y(n1647) );
  OAI21X1 U3117 ( .A(n12762), .B(n12942), .C(n1648), .Y(n5927) );
  NAND2X1 U3118 ( .A(ram[1490]), .B(n12942), .Y(n1648) );
  OAI21X1 U3119 ( .A(n12756), .B(n12942), .C(n1649), .Y(n5928) );
  NAND2X1 U3120 ( .A(ram[1491]), .B(n12942), .Y(n1649) );
  OAI21X1 U3121 ( .A(n12750), .B(n12942), .C(n1650), .Y(n5929) );
  NAND2X1 U3122 ( .A(ram[1492]), .B(n12942), .Y(n1650) );
  OAI21X1 U3123 ( .A(n12744), .B(n12942), .C(n1651), .Y(n5930) );
  NAND2X1 U3124 ( .A(ram[1493]), .B(n12942), .Y(n1651) );
  OAI21X1 U3125 ( .A(n12738), .B(n12942), .C(n1652), .Y(n5931) );
  NAND2X1 U3126 ( .A(ram[1494]), .B(n12942), .Y(n1652) );
  OAI21X1 U3127 ( .A(n12732), .B(n12942), .C(n1653), .Y(n5932) );
  NAND2X1 U3128 ( .A(ram[1495]), .B(n12942), .Y(n1653) );
  OAI21X1 U3129 ( .A(n12726), .B(n12942), .C(n1654), .Y(n5933) );
  NAND2X1 U3130 ( .A(ram[1496]), .B(n12942), .Y(n1654) );
  OAI21X1 U3131 ( .A(n12720), .B(n12942), .C(n1655), .Y(n5934) );
  NAND2X1 U3132 ( .A(ram[1497]), .B(n12942), .Y(n1655) );
  OAI21X1 U3133 ( .A(n12714), .B(n12942), .C(n1656), .Y(n5935) );
  NAND2X1 U3134 ( .A(ram[1498]), .B(n12942), .Y(n1656) );
  OAI21X1 U3135 ( .A(n12708), .B(n12942), .C(n1657), .Y(n5936) );
  NAND2X1 U3136 ( .A(ram[1499]), .B(n12942), .Y(n1657) );
  OAI21X1 U3137 ( .A(n12702), .B(n12942), .C(n1658), .Y(n5937) );
  NAND2X1 U3138 ( .A(ram[1500]), .B(n12942), .Y(n1658) );
  OAI21X1 U3139 ( .A(n12696), .B(n12942), .C(n1659), .Y(n5938) );
  NAND2X1 U3140 ( .A(ram[1501]), .B(n12942), .Y(n1659) );
  OAI21X1 U3141 ( .A(n12695), .B(n12942), .C(n1660), .Y(n5939) );
  NAND2X1 U3142 ( .A(ram[1502]), .B(n12942), .Y(n1660) );
  OAI21X1 U3143 ( .A(n12689), .B(n12942), .C(n1661), .Y(n5940) );
  NAND2X1 U3144 ( .A(ram[1503]), .B(n12942), .Y(n1661) );
  OAI21X1 U3146 ( .A(n12778), .B(n12941), .C(n1663), .Y(n5941) );
  NAND2X1 U3147 ( .A(ram[1504]), .B(n12941), .Y(n1663) );
  OAI21X1 U3148 ( .A(n12772), .B(n12941), .C(n1664), .Y(n5942) );
  NAND2X1 U3149 ( .A(ram[1505]), .B(n12941), .Y(n1664) );
  OAI21X1 U3150 ( .A(n12767), .B(n12941), .C(n1665), .Y(n5943) );
  NAND2X1 U3151 ( .A(ram[1506]), .B(n12941), .Y(n1665) );
  OAI21X1 U3152 ( .A(n12761), .B(n12941), .C(n1666), .Y(n5944) );
  NAND2X1 U3153 ( .A(ram[1507]), .B(n12941), .Y(n1666) );
  OAI21X1 U3154 ( .A(n12755), .B(n12941), .C(n1667), .Y(n5945) );
  NAND2X1 U3155 ( .A(ram[1508]), .B(n12941), .Y(n1667) );
  OAI21X1 U3156 ( .A(n12749), .B(n12941), .C(n1668), .Y(n5946) );
  NAND2X1 U3157 ( .A(ram[1509]), .B(n12941), .Y(n1668) );
  OAI21X1 U3158 ( .A(n12743), .B(n12941), .C(n1669), .Y(n5947) );
  NAND2X1 U3159 ( .A(ram[1510]), .B(n12941), .Y(n1669) );
  OAI21X1 U3160 ( .A(n12737), .B(n12941), .C(n1670), .Y(n5948) );
  NAND2X1 U3161 ( .A(ram[1511]), .B(n12941), .Y(n1670) );
  OAI21X1 U3162 ( .A(n12731), .B(n12941), .C(n1671), .Y(n5949) );
  NAND2X1 U3163 ( .A(ram[1512]), .B(n12941), .Y(n1671) );
  OAI21X1 U3164 ( .A(n12725), .B(n12941), .C(n1672), .Y(n5950) );
  NAND2X1 U3165 ( .A(ram[1513]), .B(n12941), .Y(n1672) );
  OAI21X1 U3166 ( .A(n12719), .B(n12941), .C(n1673), .Y(n5951) );
  NAND2X1 U3167 ( .A(ram[1514]), .B(n12941), .Y(n1673) );
  OAI21X1 U3168 ( .A(n12713), .B(n12941), .C(n1674), .Y(n5952) );
  NAND2X1 U3169 ( .A(ram[1515]), .B(n12941), .Y(n1674) );
  OAI21X1 U3170 ( .A(n12707), .B(n12941), .C(n1675), .Y(n5953) );
  NAND2X1 U3171 ( .A(ram[1516]), .B(n12941), .Y(n1675) );
  OAI21X1 U3172 ( .A(n12701), .B(n12941), .C(n1676), .Y(n5954) );
  NAND2X1 U3173 ( .A(ram[1517]), .B(n12941), .Y(n1676) );
  OAI21X1 U3174 ( .A(n12694), .B(n12941), .C(n1677), .Y(n5955) );
  NAND2X1 U3175 ( .A(ram[1518]), .B(n12941), .Y(n1677) );
  OAI21X1 U3176 ( .A(n12688), .B(n12941), .C(n1678), .Y(n5956) );
  NAND2X1 U3177 ( .A(ram[1519]), .B(n12941), .Y(n1678) );
  OAI21X1 U3179 ( .A(n12774), .B(n12940), .C(n1680), .Y(n5957) );
  NAND2X1 U3180 ( .A(ram[1520]), .B(n12940), .Y(n1680) );
  OAI21X1 U3181 ( .A(n12768), .B(n12940), .C(n1681), .Y(n5958) );
  NAND2X1 U3182 ( .A(ram[1521]), .B(n12940), .Y(n1681) );
  OAI21X1 U3183 ( .A(n12766), .B(n12940), .C(n1682), .Y(n5959) );
  NAND2X1 U3184 ( .A(ram[1522]), .B(n12940), .Y(n1682) );
  OAI21X1 U3185 ( .A(n12760), .B(n12940), .C(n1683), .Y(n5960) );
  NAND2X1 U3186 ( .A(ram[1523]), .B(n12940), .Y(n1683) );
  OAI21X1 U3187 ( .A(n12754), .B(n12940), .C(n1684), .Y(n5961) );
  NAND2X1 U3188 ( .A(ram[1524]), .B(n12940), .Y(n1684) );
  OAI21X1 U3189 ( .A(n12748), .B(n12940), .C(n1685), .Y(n5962) );
  NAND2X1 U3190 ( .A(ram[1525]), .B(n12940), .Y(n1685) );
  OAI21X1 U3191 ( .A(n12742), .B(n12940), .C(n1686), .Y(n5963) );
  NAND2X1 U3192 ( .A(ram[1526]), .B(n12940), .Y(n1686) );
  OAI21X1 U3193 ( .A(n12736), .B(n12940), .C(n1687), .Y(n5964) );
  NAND2X1 U3194 ( .A(ram[1527]), .B(n12940), .Y(n1687) );
  OAI21X1 U3195 ( .A(n12730), .B(n12940), .C(n1688), .Y(n5965) );
  NAND2X1 U3196 ( .A(ram[1528]), .B(n12940), .Y(n1688) );
  OAI21X1 U3197 ( .A(n12724), .B(n12940), .C(n1689), .Y(n5966) );
  NAND2X1 U3198 ( .A(ram[1529]), .B(n12940), .Y(n1689) );
  OAI21X1 U3199 ( .A(n12718), .B(n12940), .C(n1690), .Y(n5967) );
  NAND2X1 U3200 ( .A(ram[1530]), .B(n12940), .Y(n1690) );
  OAI21X1 U3201 ( .A(n12712), .B(n12940), .C(n1691), .Y(n5968) );
  NAND2X1 U3202 ( .A(ram[1531]), .B(n12940), .Y(n1691) );
  OAI21X1 U3203 ( .A(n12706), .B(n12940), .C(n1692), .Y(n5969) );
  NAND2X1 U3204 ( .A(ram[1532]), .B(n12940), .Y(n1692) );
  OAI21X1 U3205 ( .A(n12700), .B(n12940), .C(n1693), .Y(n5970) );
  NAND2X1 U3206 ( .A(ram[1533]), .B(n12940), .Y(n1693) );
  OAI21X1 U3207 ( .A(n12690), .B(n12940), .C(n1694), .Y(n5971) );
  NAND2X1 U3208 ( .A(ram[1534]), .B(n12940), .Y(n1694) );
  OAI21X1 U3209 ( .A(n12684), .B(n12940), .C(n1695), .Y(n5972) );
  NAND2X1 U3210 ( .A(ram[1535]), .B(n12940), .Y(n1695) );
  NAND3X1 U3212 ( .A(n601), .B(mem_write_en), .C(n1423), .Y(n1696) );
  OAI21X1 U3213 ( .A(n12775), .B(n12939), .C(n1698), .Y(n5973) );
  NAND2X1 U3214 ( .A(ram[1536]), .B(n12939), .Y(n1698) );
  OAI21X1 U3215 ( .A(n12769), .B(n12939), .C(n1699), .Y(n5974) );
  NAND2X1 U3216 ( .A(ram[1537]), .B(n12939), .Y(n1699) );
  OAI21X1 U3217 ( .A(n12765), .B(n12939), .C(n1700), .Y(n5975) );
  NAND2X1 U3218 ( .A(ram[1538]), .B(n12939), .Y(n1700) );
  OAI21X1 U3219 ( .A(n12759), .B(n12939), .C(n1701), .Y(n5976) );
  NAND2X1 U3220 ( .A(ram[1539]), .B(n12939), .Y(n1701) );
  OAI21X1 U3221 ( .A(n12753), .B(n12939), .C(n1702), .Y(n5977) );
  NAND2X1 U3222 ( .A(ram[1540]), .B(n12939), .Y(n1702) );
  OAI21X1 U3223 ( .A(n12747), .B(n12939), .C(n1703), .Y(n5978) );
  NAND2X1 U3224 ( .A(ram[1541]), .B(n12939), .Y(n1703) );
  OAI21X1 U3225 ( .A(n12741), .B(n12939), .C(n1704), .Y(n5979) );
  NAND2X1 U3226 ( .A(ram[1542]), .B(n12939), .Y(n1704) );
  OAI21X1 U3227 ( .A(n12735), .B(n12939), .C(n1705), .Y(n5980) );
  NAND2X1 U3228 ( .A(ram[1543]), .B(n12939), .Y(n1705) );
  OAI21X1 U3229 ( .A(n12729), .B(n12939), .C(n1706), .Y(n5981) );
  NAND2X1 U3230 ( .A(ram[1544]), .B(n12939), .Y(n1706) );
  OAI21X1 U3231 ( .A(n12723), .B(n12939), .C(n1707), .Y(n5982) );
  NAND2X1 U3232 ( .A(ram[1545]), .B(n12939), .Y(n1707) );
  OAI21X1 U3233 ( .A(n12717), .B(n12939), .C(n1708), .Y(n5983) );
  NAND2X1 U3234 ( .A(ram[1546]), .B(n12939), .Y(n1708) );
  OAI21X1 U3235 ( .A(n12711), .B(n12939), .C(n1709), .Y(n5984) );
  NAND2X1 U3236 ( .A(ram[1547]), .B(n12939), .Y(n1709) );
  OAI21X1 U3237 ( .A(n12705), .B(n12939), .C(n1710), .Y(n5985) );
  NAND2X1 U3238 ( .A(ram[1548]), .B(n12939), .Y(n1710) );
  OAI21X1 U3239 ( .A(n12699), .B(n12939), .C(n1711), .Y(n5986) );
  NAND2X1 U3240 ( .A(ram[1549]), .B(n12939), .Y(n1711) );
  OAI21X1 U3241 ( .A(n12691), .B(n12939), .C(n1712), .Y(n5987) );
  NAND2X1 U3242 ( .A(ram[1550]), .B(n12939), .Y(n1712) );
  OAI21X1 U3243 ( .A(n12685), .B(n12939), .C(n1713), .Y(n5988) );
  NAND2X1 U3244 ( .A(ram[1551]), .B(n12939), .Y(n1713) );
  OAI21X1 U3246 ( .A(n12778), .B(n12938), .C(n1715), .Y(n5989) );
  NAND2X1 U3247 ( .A(ram[1552]), .B(n12938), .Y(n1715) );
  OAI21X1 U3248 ( .A(n12772), .B(n12938), .C(n1716), .Y(n5990) );
  NAND2X1 U3249 ( .A(ram[1553]), .B(n12938), .Y(n1716) );
  OAI21X1 U3250 ( .A(n12763), .B(n12938), .C(n1717), .Y(n5991) );
  NAND2X1 U3251 ( .A(ram[1554]), .B(n12938), .Y(n1717) );
  OAI21X1 U3252 ( .A(n12757), .B(n12938), .C(n1718), .Y(n5992) );
  NAND2X1 U3253 ( .A(ram[1555]), .B(n12938), .Y(n1718) );
  OAI21X1 U3254 ( .A(n12751), .B(n12938), .C(n1719), .Y(n5993) );
  NAND2X1 U3255 ( .A(ram[1556]), .B(n12938), .Y(n1719) );
  OAI21X1 U3256 ( .A(n12745), .B(n12938), .C(n1720), .Y(n5994) );
  NAND2X1 U3257 ( .A(ram[1557]), .B(n12938), .Y(n1720) );
  OAI21X1 U3258 ( .A(n12739), .B(n12938), .C(n1721), .Y(n5995) );
  NAND2X1 U3259 ( .A(ram[1558]), .B(n12938), .Y(n1721) );
  OAI21X1 U3260 ( .A(n12733), .B(n12938), .C(n1722), .Y(n5996) );
  NAND2X1 U3261 ( .A(ram[1559]), .B(n12938), .Y(n1722) );
  OAI21X1 U3262 ( .A(n12727), .B(n12938), .C(n1723), .Y(n5997) );
  NAND2X1 U3263 ( .A(ram[1560]), .B(n12938), .Y(n1723) );
  OAI21X1 U3264 ( .A(n12721), .B(n12938), .C(n1724), .Y(n5998) );
  NAND2X1 U3265 ( .A(ram[1561]), .B(n12938), .Y(n1724) );
  OAI21X1 U3266 ( .A(n12715), .B(n12938), .C(n1725), .Y(n5999) );
  NAND2X1 U3267 ( .A(ram[1562]), .B(n12938), .Y(n1725) );
  OAI21X1 U3268 ( .A(n12709), .B(n12938), .C(n1726), .Y(n6000) );
  NAND2X1 U3269 ( .A(ram[1563]), .B(n12938), .Y(n1726) );
  OAI21X1 U3270 ( .A(n12703), .B(n12938), .C(n1727), .Y(n6001) );
  NAND2X1 U3271 ( .A(ram[1564]), .B(n12938), .Y(n1727) );
  OAI21X1 U3272 ( .A(n12697), .B(n12938), .C(n1728), .Y(n6002) );
  NAND2X1 U3273 ( .A(ram[1565]), .B(n12938), .Y(n1728) );
  OAI21X1 U3274 ( .A(n12694), .B(n12938), .C(n1729), .Y(n6003) );
  NAND2X1 U3275 ( .A(ram[1566]), .B(n12938), .Y(n1729) );
  OAI21X1 U3276 ( .A(n12688), .B(n12938), .C(n1730), .Y(n6004) );
  NAND2X1 U3277 ( .A(ram[1567]), .B(n12938), .Y(n1730) );
  OAI21X1 U3279 ( .A(n12777), .B(n12937), .C(n1732), .Y(n6005) );
  NAND2X1 U3280 ( .A(ram[1568]), .B(n12937), .Y(n1732) );
  OAI21X1 U3281 ( .A(n12771), .B(n12937), .C(n1733), .Y(n6006) );
  NAND2X1 U3282 ( .A(ram[1569]), .B(n12937), .Y(n1733) );
  OAI21X1 U3283 ( .A(n12766), .B(n12937), .C(n1734), .Y(n6007) );
  NAND2X1 U3284 ( .A(ram[1570]), .B(n12937), .Y(n1734) );
  OAI21X1 U3285 ( .A(n12760), .B(n12937), .C(n1735), .Y(n6008) );
  NAND2X1 U3286 ( .A(ram[1571]), .B(n12937), .Y(n1735) );
  OAI21X1 U3287 ( .A(n12754), .B(n12937), .C(n1736), .Y(n6009) );
  NAND2X1 U3288 ( .A(ram[1572]), .B(n12937), .Y(n1736) );
  OAI21X1 U3289 ( .A(n12748), .B(n12937), .C(n1737), .Y(n6010) );
  NAND2X1 U3290 ( .A(ram[1573]), .B(n12937), .Y(n1737) );
  OAI21X1 U3291 ( .A(n12742), .B(n12937), .C(n1738), .Y(n6011) );
  NAND2X1 U3292 ( .A(ram[1574]), .B(n12937), .Y(n1738) );
  OAI21X1 U3293 ( .A(n12736), .B(n12937), .C(n1739), .Y(n6012) );
  NAND2X1 U3294 ( .A(ram[1575]), .B(n12937), .Y(n1739) );
  OAI21X1 U3295 ( .A(n12730), .B(n12937), .C(n1740), .Y(n6013) );
  NAND2X1 U3296 ( .A(ram[1576]), .B(n12937), .Y(n1740) );
  OAI21X1 U3297 ( .A(n12724), .B(n12937), .C(n1741), .Y(n6014) );
  NAND2X1 U3298 ( .A(ram[1577]), .B(n12937), .Y(n1741) );
  OAI21X1 U3299 ( .A(n12718), .B(n12937), .C(n1742), .Y(n6015) );
  NAND2X1 U3300 ( .A(ram[1578]), .B(n12937), .Y(n1742) );
  OAI21X1 U3301 ( .A(n12712), .B(n12937), .C(n1743), .Y(n6016) );
  NAND2X1 U3302 ( .A(ram[1579]), .B(n12937), .Y(n1743) );
  OAI21X1 U3303 ( .A(n12706), .B(n12937), .C(n1744), .Y(n6017) );
  NAND2X1 U3304 ( .A(ram[1580]), .B(n12937), .Y(n1744) );
  OAI21X1 U3305 ( .A(n12700), .B(n12937), .C(n1745), .Y(n6018) );
  NAND2X1 U3306 ( .A(ram[1581]), .B(n12937), .Y(n1745) );
  OAI21X1 U3307 ( .A(n12693), .B(n12937), .C(n1746), .Y(n6019) );
  NAND2X1 U3308 ( .A(ram[1582]), .B(n12937), .Y(n1746) );
  OAI21X1 U3309 ( .A(n12687), .B(n12937), .C(n1747), .Y(n6020) );
  NAND2X1 U3310 ( .A(ram[1583]), .B(n12937), .Y(n1747) );
  OAI21X1 U3312 ( .A(n12774), .B(n12936), .C(n1749), .Y(n6021) );
  NAND2X1 U3313 ( .A(ram[1584]), .B(n12936), .Y(n1749) );
  OAI21X1 U3314 ( .A(n12768), .B(n12936), .C(n1750), .Y(n6022) );
  NAND2X1 U3315 ( .A(ram[1585]), .B(n12936), .Y(n1750) );
  OAI21X1 U3316 ( .A(n12764), .B(n12936), .C(n1751), .Y(n6023) );
  NAND2X1 U3317 ( .A(ram[1586]), .B(n12936), .Y(n1751) );
  OAI21X1 U3318 ( .A(n12758), .B(n12936), .C(n1752), .Y(n6024) );
  NAND2X1 U3319 ( .A(ram[1587]), .B(n12936), .Y(n1752) );
  OAI21X1 U3320 ( .A(n12752), .B(n12936), .C(n1753), .Y(n6025) );
  NAND2X1 U3321 ( .A(ram[1588]), .B(n12936), .Y(n1753) );
  OAI21X1 U3322 ( .A(n12746), .B(n12936), .C(n1754), .Y(n6026) );
  NAND2X1 U3323 ( .A(ram[1589]), .B(n12936), .Y(n1754) );
  OAI21X1 U3324 ( .A(n12740), .B(n12936), .C(n1755), .Y(n6027) );
  NAND2X1 U3325 ( .A(ram[1590]), .B(n12936), .Y(n1755) );
  OAI21X1 U3326 ( .A(n12734), .B(n12936), .C(n1756), .Y(n6028) );
  NAND2X1 U3327 ( .A(ram[1591]), .B(n12936), .Y(n1756) );
  OAI21X1 U3328 ( .A(n12728), .B(n12936), .C(n1757), .Y(n6029) );
  NAND2X1 U3329 ( .A(ram[1592]), .B(n12936), .Y(n1757) );
  OAI21X1 U3330 ( .A(n12722), .B(n12936), .C(n1758), .Y(n6030) );
  NAND2X1 U3331 ( .A(ram[1593]), .B(n12936), .Y(n1758) );
  OAI21X1 U3332 ( .A(n12716), .B(n12936), .C(n1759), .Y(n6031) );
  NAND2X1 U3333 ( .A(ram[1594]), .B(n12936), .Y(n1759) );
  OAI21X1 U3334 ( .A(n12710), .B(n12936), .C(n1760), .Y(n6032) );
  NAND2X1 U3335 ( .A(ram[1595]), .B(n12936), .Y(n1760) );
  OAI21X1 U3336 ( .A(n12704), .B(n12936), .C(n1761), .Y(n6033) );
  NAND2X1 U3337 ( .A(ram[1596]), .B(n12936), .Y(n1761) );
  OAI21X1 U3338 ( .A(n12698), .B(n12936), .C(n1762), .Y(n6034) );
  NAND2X1 U3339 ( .A(ram[1597]), .B(n12936), .Y(n1762) );
  OAI21X1 U3340 ( .A(n12690), .B(n12936), .C(n1763), .Y(n6035) );
  NAND2X1 U3341 ( .A(ram[1598]), .B(n12936), .Y(n1763) );
  OAI21X1 U3342 ( .A(n12684), .B(n12936), .C(n1764), .Y(n6036) );
  NAND2X1 U3343 ( .A(ram[1599]), .B(n12936), .Y(n1764) );
  OAI21X1 U3345 ( .A(n12775), .B(n12935), .C(n1766), .Y(n6037) );
  NAND2X1 U3346 ( .A(ram[1600]), .B(n12935), .Y(n1766) );
  OAI21X1 U3347 ( .A(n12769), .B(n12935), .C(n1767), .Y(n6038) );
  NAND2X1 U3348 ( .A(ram[1601]), .B(n12935), .Y(n1767) );
  OAI21X1 U3349 ( .A(n12765), .B(n12935), .C(n1768), .Y(n6039) );
  NAND2X1 U3350 ( .A(ram[1602]), .B(n12935), .Y(n1768) );
  OAI21X1 U3351 ( .A(n12759), .B(n12935), .C(n1769), .Y(n6040) );
  NAND2X1 U3352 ( .A(ram[1603]), .B(n12935), .Y(n1769) );
  OAI21X1 U3353 ( .A(n12753), .B(n12935), .C(n1770), .Y(n6041) );
  NAND2X1 U3354 ( .A(ram[1604]), .B(n12935), .Y(n1770) );
  OAI21X1 U3355 ( .A(n12747), .B(n12935), .C(n1771), .Y(n6042) );
  NAND2X1 U3356 ( .A(ram[1605]), .B(n12935), .Y(n1771) );
  OAI21X1 U3357 ( .A(n12741), .B(n12935), .C(n1772), .Y(n6043) );
  NAND2X1 U3358 ( .A(ram[1606]), .B(n12935), .Y(n1772) );
  OAI21X1 U3359 ( .A(n12735), .B(n12935), .C(n1773), .Y(n6044) );
  NAND2X1 U3360 ( .A(ram[1607]), .B(n12935), .Y(n1773) );
  OAI21X1 U3361 ( .A(n12729), .B(n12935), .C(n1774), .Y(n6045) );
  NAND2X1 U3362 ( .A(ram[1608]), .B(n12935), .Y(n1774) );
  OAI21X1 U3363 ( .A(n12723), .B(n12935), .C(n1775), .Y(n6046) );
  NAND2X1 U3364 ( .A(ram[1609]), .B(n12935), .Y(n1775) );
  OAI21X1 U3365 ( .A(n12717), .B(n12935), .C(n1776), .Y(n6047) );
  NAND2X1 U3366 ( .A(ram[1610]), .B(n12935), .Y(n1776) );
  OAI21X1 U3367 ( .A(n12711), .B(n12935), .C(n1777), .Y(n6048) );
  NAND2X1 U3368 ( .A(ram[1611]), .B(n12935), .Y(n1777) );
  OAI21X1 U3369 ( .A(n12705), .B(n12935), .C(n1778), .Y(n6049) );
  NAND2X1 U3370 ( .A(ram[1612]), .B(n12935), .Y(n1778) );
  OAI21X1 U3371 ( .A(n12699), .B(n12935), .C(n1779), .Y(n6050) );
  NAND2X1 U3372 ( .A(ram[1613]), .B(n12935), .Y(n1779) );
  OAI21X1 U3373 ( .A(n12691), .B(n12935), .C(n1780), .Y(n6051) );
  NAND2X1 U3374 ( .A(ram[1614]), .B(n12935), .Y(n1780) );
  OAI21X1 U3375 ( .A(n12685), .B(n12935), .C(n1781), .Y(n6052) );
  NAND2X1 U3376 ( .A(ram[1615]), .B(n12935), .Y(n1781) );
  OAI21X1 U3378 ( .A(n12777), .B(n12934), .C(n1783), .Y(n6053) );
  NAND2X1 U3379 ( .A(ram[1616]), .B(n12934), .Y(n1783) );
  OAI21X1 U3380 ( .A(n12771), .B(n12934), .C(n1784), .Y(n6054) );
  NAND2X1 U3381 ( .A(ram[1617]), .B(n12934), .Y(n1784) );
  OAI21X1 U3382 ( .A(n12764), .B(n12934), .C(n1785), .Y(n6055) );
  NAND2X1 U3383 ( .A(ram[1618]), .B(n12934), .Y(n1785) );
  OAI21X1 U3384 ( .A(n12758), .B(n12934), .C(n1786), .Y(n6056) );
  NAND2X1 U3385 ( .A(ram[1619]), .B(n12934), .Y(n1786) );
  OAI21X1 U3386 ( .A(n12752), .B(n12934), .C(n1787), .Y(n6057) );
  NAND2X1 U3387 ( .A(ram[1620]), .B(n12934), .Y(n1787) );
  OAI21X1 U3388 ( .A(n12746), .B(n12934), .C(n1788), .Y(n6058) );
  NAND2X1 U3389 ( .A(ram[1621]), .B(n12934), .Y(n1788) );
  OAI21X1 U3390 ( .A(n12740), .B(n12934), .C(n1789), .Y(n6059) );
  NAND2X1 U3391 ( .A(ram[1622]), .B(n12934), .Y(n1789) );
  OAI21X1 U3392 ( .A(n12734), .B(n12934), .C(n1790), .Y(n6060) );
  NAND2X1 U3393 ( .A(ram[1623]), .B(n12934), .Y(n1790) );
  OAI21X1 U3394 ( .A(n12728), .B(n12934), .C(n1791), .Y(n6061) );
  NAND2X1 U3395 ( .A(ram[1624]), .B(n12934), .Y(n1791) );
  OAI21X1 U3396 ( .A(n12722), .B(n12934), .C(n1792), .Y(n6062) );
  NAND2X1 U3397 ( .A(ram[1625]), .B(n12934), .Y(n1792) );
  OAI21X1 U3398 ( .A(n12716), .B(n12934), .C(n1793), .Y(n6063) );
  NAND2X1 U3399 ( .A(ram[1626]), .B(n12934), .Y(n1793) );
  OAI21X1 U3400 ( .A(n12710), .B(n12934), .C(n1794), .Y(n6064) );
  NAND2X1 U3401 ( .A(ram[1627]), .B(n12934), .Y(n1794) );
  OAI21X1 U3402 ( .A(n12704), .B(n12934), .C(n1795), .Y(n6065) );
  NAND2X1 U3403 ( .A(ram[1628]), .B(n12934), .Y(n1795) );
  OAI21X1 U3404 ( .A(n12698), .B(n12934), .C(n1796), .Y(n6066) );
  NAND2X1 U3405 ( .A(ram[1629]), .B(n12934), .Y(n1796) );
  OAI21X1 U3406 ( .A(n12693), .B(n12934), .C(n1797), .Y(n6067) );
  NAND2X1 U3407 ( .A(ram[1630]), .B(n12934), .Y(n1797) );
  OAI21X1 U3408 ( .A(n12687), .B(n12934), .C(n1798), .Y(n6068) );
  NAND2X1 U3409 ( .A(ram[1631]), .B(n12934), .Y(n1798) );
  OAI21X1 U3411 ( .A(n12778), .B(n12933), .C(n1800), .Y(n6069) );
  NAND2X1 U3412 ( .A(ram[1632]), .B(n12933), .Y(n1800) );
  OAI21X1 U3413 ( .A(n12772), .B(n12933), .C(n1801), .Y(n6070) );
  NAND2X1 U3414 ( .A(ram[1633]), .B(n12933), .Y(n1801) );
  OAI21X1 U3415 ( .A(n12765), .B(n12933), .C(n1802), .Y(n6071) );
  NAND2X1 U3416 ( .A(ram[1634]), .B(n12933), .Y(n1802) );
  OAI21X1 U3417 ( .A(n12759), .B(n12933), .C(n1803), .Y(n6072) );
  NAND2X1 U3418 ( .A(ram[1635]), .B(n12933), .Y(n1803) );
  OAI21X1 U3419 ( .A(n12753), .B(n12933), .C(n1804), .Y(n6073) );
  NAND2X1 U3420 ( .A(ram[1636]), .B(n12933), .Y(n1804) );
  OAI21X1 U3421 ( .A(n12747), .B(n12933), .C(n1805), .Y(n6074) );
  NAND2X1 U3422 ( .A(ram[1637]), .B(n12933), .Y(n1805) );
  OAI21X1 U3423 ( .A(n12741), .B(n12933), .C(n1806), .Y(n6075) );
  NAND2X1 U3424 ( .A(ram[1638]), .B(n12933), .Y(n1806) );
  OAI21X1 U3425 ( .A(n12735), .B(n12933), .C(n1807), .Y(n6076) );
  NAND2X1 U3426 ( .A(ram[1639]), .B(n12933), .Y(n1807) );
  OAI21X1 U3427 ( .A(n12729), .B(n12933), .C(n1808), .Y(n6077) );
  NAND2X1 U3428 ( .A(ram[1640]), .B(n12933), .Y(n1808) );
  OAI21X1 U3429 ( .A(n12723), .B(n12933), .C(n1809), .Y(n6078) );
  NAND2X1 U3430 ( .A(ram[1641]), .B(n12933), .Y(n1809) );
  OAI21X1 U3431 ( .A(n12717), .B(n12933), .C(n1810), .Y(n6079) );
  NAND2X1 U3432 ( .A(ram[1642]), .B(n12933), .Y(n1810) );
  OAI21X1 U3433 ( .A(n12711), .B(n12933), .C(n1811), .Y(n6080) );
  NAND2X1 U3434 ( .A(ram[1643]), .B(n12933), .Y(n1811) );
  OAI21X1 U3435 ( .A(n12705), .B(n12933), .C(n1812), .Y(n6081) );
  NAND2X1 U3436 ( .A(ram[1644]), .B(n12933), .Y(n1812) );
  OAI21X1 U3437 ( .A(n12699), .B(n12933), .C(n1813), .Y(n6082) );
  NAND2X1 U3438 ( .A(ram[1645]), .B(n12933), .Y(n1813) );
  OAI21X1 U3439 ( .A(n12694), .B(n12933), .C(n1814), .Y(n6083) );
  NAND2X1 U3440 ( .A(ram[1646]), .B(n12933), .Y(n1814) );
  OAI21X1 U3441 ( .A(n12688), .B(n12933), .C(n1815), .Y(n6084) );
  NAND2X1 U3442 ( .A(ram[1647]), .B(n12933), .Y(n1815) );
  OAI21X1 U3444 ( .A(n12774), .B(n12932), .C(n1817), .Y(n6085) );
  NAND2X1 U3445 ( .A(ram[1648]), .B(n12932), .Y(n1817) );
  OAI21X1 U3446 ( .A(n12768), .B(n12932), .C(n1818), .Y(n6086) );
  NAND2X1 U3447 ( .A(ram[1649]), .B(n12932), .Y(n1818) );
  OAI21X1 U3448 ( .A(n12765), .B(n12932), .C(n1819), .Y(n6087) );
  NAND2X1 U3449 ( .A(ram[1650]), .B(n12932), .Y(n1819) );
  OAI21X1 U3450 ( .A(n12759), .B(n12932), .C(n1820), .Y(n6088) );
  NAND2X1 U3451 ( .A(ram[1651]), .B(n12932), .Y(n1820) );
  OAI21X1 U3452 ( .A(n12753), .B(n12932), .C(n1821), .Y(n6089) );
  NAND2X1 U3453 ( .A(ram[1652]), .B(n12932), .Y(n1821) );
  OAI21X1 U3454 ( .A(n12747), .B(n12932), .C(n1822), .Y(n6090) );
  NAND2X1 U3455 ( .A(ram[1653]), .B(n12932), .Y(n1822) );
  OAI21X1 U3456 ( .A(n12741), .B(n12932), .C(n1823), .Y(n6091) );
  NAND2X1 U3457 ( .A(ram[1654]), .B(n12932), .Y(n1823) );
  OAI21X1 U3458 ( .A(n12735), .B(n12932), .C(n1824), .Y(n6092) );
  NAND2X1 U3459 ( .A(ram[1655]), .B(n12932), .Y(n1824) );
  OAI21X1 U3460 ( .A(n12729), .B(n12932), .C(n1825), .Y(n6093) );
  NAND2X1 U3461 ( .A(ram[1656]), .B(n12932), .Y(n1825) );
  OAI21X1 U3462 ( .A(n12723), .B(n12932), .C(n1826), .Y(n6094) );
  NAND2X1 U3463 ( .A(ram[1657]), .B(n12932), .Y(n1826) );
  OAI21X1 U3464 ( .A(n12717), .B(n12932), .C(n1827), .Y(n6095) );
  NAND2X1 U3465 ( .A(ram[1658]), .B(n12932), .Y(n1827) );
  OAI21X1 U3466 ( .A(n12711), .B(n12932), .C(n1828), .Y(n6096) );
  NAND2X1 U3467 ( .A(ram[1659]), .B(n12932), .Y(n1828) );
  OAI21X1 U3468 ( .A(n12705), .B(n12932), .C(n1829), .Y(n6097) );
  NAND2X1 U3469 ( .A(ram[1660]), .B(n12932), .Y(n1829) );
  OAI21X1 U3470 ( .A(n12699), .B(n12932), .C(n1830), .Y(n6098) );
  NAND2X1 U3471 ( .A(ram[1661]), .B(n12932), .Y(n1830) );
  OAI21X1 U3472 ( .A(n12690), .B(n12932), .C(n1831), .Y(n6099) );
  NAND2X1 U3473 ( .A(ram[1662]), .B(n12932), .Y(n1831) );
  OAI21X1 U3474 ( .A(n12684), .B(n12932), .C(n1832), .Y(n6100) );
  NAND2X1 U3475 ( .A(ram[1663]), .B(n12932), .Y(n1832) );
  OAI21X1 U3477 ( .A(n12776), .B(n12931), .C(n1834), .Y(n6101) );
  NAND2X1 U3478 ( .A(ram[1664]), .B(n12931), .Y(n1834) );
  OAI21X1 U3479 ( .A(n12770), .B(n12931), .C(n1835), .Y(n6102) );
  NAND2X1 U3480 ( .A(ram[1665]), .B(n12931), .Y(n1835) );
  OAI21X1 U3481 ( .A(n12767), .B(n12931), .C(n1836), .Y(n6103) );
  NAND2X1 U3482 ( .A(ram[1666]), .B(n12931), .Y(n1836) );
  OAI21X1 U3483 ( .A(n12761), .B(n12931), .C(n1837), .Y(n6104) );
  NAND2X1 U3484 ( .A(ram[1667]), .B(n12931), .Y(n1837) );
  OAI21X1 U3485 ( .A(n12755), .B(n12931), .C(n1838), .Y(n6105) );
  NAND2X1 U3486 ( .A(ram[1668]), .B(n12931), .Y(n1838) );
  OAI21X1 U3487 ( .A(n12749), .B(n12931), .C(n1839), .Y(n6106) );
  NAND2X1 U3488 ( .A(ram[1669]), .B(n12931), .Y(n1839) );
  OAI21X1 U3489 ( .A(n12743), .B(n12931), .C(n1840), .Y(n6107) );
  NAND2X1 U3490 ( .A(ram[1670]), .B(n12931), .Y(n1840) );
  OAI21X1 U3491 ( .A(n12737), .B(n12931), .C(n1841), .Y(n6108) );
  NAND2X1 U3492 ( .A(ram[1671]), .B(n12931), .Y(n1841) );
  OAI21X1 U3493 ( .A(n12731), .B(n12931), .C(n1842), .Y(n6109) );
  NAND2X1 U3494 ( .A(ram[1672]), .B(n12931), .Y(n1842) );
  OAI21X1 U3495 ( .A(n12725), .B(n12931), .C(n1843), .Y(n6110) );
  NAND2X1 U3496 ( .A(ram[1673]), .B(n12931), .Y(n1843) );
  OAI21X1 U3497 ( .A(n12719), .B(n12931), .C(n1844), .Y(n6111) );
  NAND2X1 U3498 ( .A(ram[1674]), .B(n12931), .Y(n1844) );
  OAI21X1 U3499 ( .A(n12713), .B(n12931), .C(n1845), .Y(n6112) );
  NAND2X1 U3500 ( .A(ram[1675]), .B(n12931), .Y(n1845) );
  OAI21X1 U3501 ( .A(n12707), .B(n12931), .C(n1846), .Y(n6113) );
  NAND2X1 U3502 ( .A(ram[1676]), .B(n12931), .Y(n1846) );
  OAI21X1 U3503 ( .A(n12701), .B(n12931), .C(n1847), .Y(n6114) );
  NAND2X1 U3504 ( .A(ram[1677]), .B(n12931), .Y(n1847) );
  OAI21X1 U3505 ( .A(n12692), .B(n12931), .C(n1848), .Y(n6115) );
  NAND2X1 U3506 ( .A(ram[1678]), .B(n12931), .Y(n1848) );
  OAI21X1 U3507 ( .A(n12686), .B(n12931), .C(n1849), .Y(n6116) );
  NAND2X1 U3508 ( .A(ram[1679]), .B(n12931), .Y(n1849) );
  OAI21X1 U3510 ( .A(n12775), .B(n12930), .C(n1851), .Y(n6117) );
  NAND2X1 U3511 ( .A(ram[1680]), .B(n12930), .Y(n1851) );
  OAI21X1 U3512 ( .A(n12769), .B(n12930), .C(n1852), .Y(n6118) );
  NAND2X1 U3513 ( .A(ram[1681]), .B(n12930), .Y(n1852) );
  OAI21X1 U3514 ( .A(n12766), .B(n12930), .C(n1853), .Y(n6119) );
  NAND2X1 U3515 ( .A(ram[1682]), .B(n12930), .Y(n1853) );
  OAI21X1 U3516 ( .A(n12760), .B(n12930), .C(n1854), .Y(n6120) );
  NAND2X1 U3517 ( .A(ram[1683]), .B(n12930), .Y(n1854) );
  OAI21X1 U3518 ( .A(n12754), .B(n12930), .C(n1855), .Y(n6121) );
  NAND2X1 U3519 ( .A(ram[1684]), .B(n12930), .Y(n1855) );
  OAI21X1 U3520 ( .A(n12748), .B(n12930), .C(n1856), .Y(n6122) );
  NAND2X1 U3521 ( .A(ram[1685]), .B(n12930), .Y(n1856) );
  OAI21X1 U3522 ( .A(n12742), .B(n12930), .C(n1857), .Y(n6123) );
  NAND2X1 U3523 ( .A(ram[1686]), .B(n12930), .Y(n1857) );
  OAI21X1 U3524 ( .A(n12736), .B(n12930), .C(n1858), .Y(n6124) );
  NAND2X1 U3525 ( .A(ram[1687]), .B(n12930), .Y(n1858) );
  OAI21X1 U3526 ( .A(n12730), .B(n12930), .C(n1859), .Y(n6125) );
  NAND2X1 U3527 ( .A(ram[1688]), .B(n12930), .Y(n1859) );
  OAI21X1 U3528 ( .A(n12724), .B(n12930), .C(n1860), .Y(n6126) );
  NAND2X1 U3529 ( .A(ram[1689]), .B(n12930), .Y(n1860) );
  OAI21X1 U3530 ( .A(n12718), .B(n12930), .C(n1861), .Y(n6127) );
  NAND2X1 U3531 ( .A(ram[1690]), .B(n12930), .Y(n1861) );
  OAI21X1 U3532 ( .A(n12712), .B(n12930), .C(n1862), .Y(n6128) );
  NAND2X1 U3533 ( .A(ram[1691]), .B(n12930), .Y(n1862) );
  OAI21X1 U3534 ( .A(n12706), .B(n12930), .C(n1863), .Y(n6129) );
  NAND2X1 U3535 ( .A(ram[1692]), .B(n12930), .Y(n1863) );
  OAI21X1 U3536 ( .A(n12700), .B(n12930), .C(n1864), .Y(n6130) );
  NAND2X1 U3537 ( .A(ram[1693]), .B(n12930), .Y(n1864) );
  OAI21X1 U3538 ( .A(n12691), .B(n12930), .C(n1865), .Y(n6131) );
  NAND2X1 U3539 ( .A(ram[1694]), .B(n12930), .Y(n1865) );
  OAI21X1 U3540 ( .A(n12685), .B(n12930), .C(n1866), .Y(n6132) );
  NAND2X1 U3541 ( .A(ram[1695]), .B(n12930), .Y(n1866) );
  OAI21X1 U3543 ( .A(n12774), .B(n12929), .C(n1868), .Y(n6133) );
  NAND2X1 U3544 ( .A(ram[1696]), .B(n12929), .Y(n1868) );
  OAI21X1 U3545 ( .A(n12768), .B(n12929), .C(n1869), .Y(n6134) );
  NAND2X1 U3546 ( .A(ram[1697]), .B(n12929), .Y(n1869) );
  OAI21X1 U3547 ( .A(n12765), .B(n12929), .C(n1870), .Y(n6135) );
  NAND2X1 U3548 ( .A(ram[1698]), .B(n12929), .Y(n1870) );
  OAI21X1 U3549 ( .A(n12759), .B(n12929), .C(n1871), .Y(n6136) );
  NAND2X1 U3550 ( .A(ram[1699]), .B(n12929), .Y(n1871) );
  OAI21X1 U3551 ( .A(n12753), .B(n12929), .C(n1872), .Y(n6137) );
  NAND2X1 U3552 ( .A(ram[1700]), .B(n12929), .Y(n1872) );
  OAI21X1 U3553 ( .A(n12747), .B(n12929), .C(n1873), .Y(n6138) );
  NAND2X1 U3554 ( .A(ram[1701]), .B(n12929), .Y(n1873) );
  OAI21X1 U3555 ( .A(n12741), .B(n12929), .C(n1874), .Y(n6139) );
  NAND2X1 U3556 ( .A(ram[1702]), .B(n12929), .Y(n1874) );
  OAI21X1 U3557 ( .A(n12735), .B(n12929), .C(n1875), .Y(n6140) );
  NAND2X1 U3558 ( .A(ram[1703]), .B(n12929), .Y(n1875) );
  OAI21X1 U3559 ( .A(n12729), .B(n12929), .C(n1876), .Y(n6141) );
  NAND2X1 U3560 ( .A(ram[1704]), .B(n12929), .Y(n1876) );
  OAI21X1 U3561 ( .A(n12723), .B(n12929), .C(n1877), .Y(n6142) );
  NAND2X1 U3562 ( .A(ram[1705]), .B(n12929), .Y(n1877) );
  OAI21X1 U3563 ( .A(n12717), .B(n12929), .C(n1878), .Y(n6143) );
  NAND2X1 U3564 ( .A(ram[1706]), .B(n12929), .Y(n1878) );
  OAI21X1 U3565 ( .A(n12711), .B(n12929), .C(n1879), .Y(n6144) );
  NAND2X1 U3566 ( .A(ram[1707]), .B(n12929), .Y(n1879) );
  OAI21X1 U3567 ( .A(n12705), .B(n12929), .C(n1880), .Y(n6145) );
  NAND2X1 U3568 ( .A(ram[1708]), .B(n12929), .Y(n1880) );
  OAI21X1 U3569 ( .A(n12699), .B(n12929), .C(n1881), .Y(n6146) );
  NAND2X1 U3570 ( .A(ram[1709]), .B(n12929), .Y(n1881) );
  OAI21X1 U3571 ( .A(n12690), .B(n12929), .C(n1882), .Y(n6147) );
  NAND2X1 U3572 ( .A(ram[1710]), .B(n12929), .Y(n1882) );
  OAI21X1 U3573 ( .A(n12684), .B(n12929), .C(n1883), .Y(n6148) );
  NAND2X1 U3574 ( .A(ram[1711]), .B(n12929), .Y(n1883) );
  OAI21X1 U3576 ( .A(n12779), .B(n12928), .C(n1885), .Y(n6149) );
  NAND2X1 U3577 ( .A(ram[1712]), .B(n12928), .Y(n1885) );
  OAI21X1 U3578 ( .A(n12773), .B(n12928), .C(n1886), .Y(n6150) );
  NAND2X1 U3579 ( .A(ram[1713]), .B(n12928), .Y(n1886) );
  OAI21X1 U3580 ( .A(n12767), .B(n12928), .C(n1887), .Y(n6151) );
  NAND2X1 U3581 ( .A(ram[1714]), .B(n12928), .Y(n1887) );
  OAI21X1 U3582 ( .A(n12761), .B(n12928), .C(n1888), .Y(n6152) );
  NAND2X1 U3583 ( .A(ram[1715]), .B(n12928), .Y(n1888) );
  OAI21X1 U3584 ( .A(n12755), .B(n12928), .C(n1889), .Y(n6153) );
  NAND2X1 U3585 ( .A(ram[1716]), .B(n12928), .Y(n1889) );
  OAI21X1 U3586 ( .A(n12749), .B(n12928), .C(n1890), .Y(n6154) );
  NAND2X1 U3587 ( .A(ram[1717]), .B(n12928), .Y(n1890) );
  OAI21X1 U3588 ( .A(n12743), .B(n12928), .C(n1891), .Y(n6155) );
  NAND2X1 U3589 ( .A(ram[1718]), .B(n12928), .Y(n1891) );
  OAI21X1 U3590 ( .A(n12737), .B(n12928), .C(n1892), .Y(n6156) );
  NAND2X1 U3591 ( .A(ram[1719]), .B(n12928), .Y(n1892) );
  OAI21X1 U3592 ( .A(n12731), .B(n12928), .C(n1893), .Y(n6157) );
  NAND2X1 U3593 ( .A(ram[1720]), .B(n12928), .Y(n1893) );
  OAI21X1 U3594 ( .A(n12725), .B(n12928), .C(n1894), .Y(n6158) );
  NAND2X1 U3595 ( .A(ram[1721]), .B(n12928), .Y(n1894) );
  OAI21X1 U3596 ( .A(n12719), .B(n12928), .C(n1895), .Y(n6159) );
  NAND2X1 U3597 ( .A(ram[1722]), .B(n12928), .Y(n1895) );
  OAI21X1 U3598 ( .A(n12713), .B(n12928), .C(n1896), .Y(n6160) );
  NAND2X1 U3599 ( .A(ram[1723]), .B(n12928), .Y(n1896) );
  OAI21X1 U3600 ( .A(n12707), .B(n12928), .C(n1897), .Y(n6161) );
  NAND2X1 U3601 ( .A(ram[1724]), .B(n12928), .Y(n1897) );
  OAI21X1 U3602 ( .A(n12701), .B(n12928), .C(n1898), .Y(n6162) );
  NAND2X1 U3603 ( .A(ram[1725]), .B(n12928), .Y(n1898) );
  OAI21X1 U3604 ( .A(n12695), .B(n12928), .C(n1899), .Y(n6163) );
  NAND2X1 U3605 ( .A(ram[1726]), .B(n12928), .Y(n1899) );
  OAI21X1 U3606 ( .A(n12689), .B(n12928), .C(n1900), .Y(n6164) );
  NAND2X1 U3607 ( .A(ram[1727]), .B(n12928), .Y(n1900) );
  OAI21X1 U3609 ( .A(n12778), .B(n12927), .C(n1902), .Y(n6165) );
  NAND2X1 U3610 ( .A(ram[1728]), .B(n12927), .Y(n1902) );
  OAI21X1 U3611 ( .A(n12772), .B(n12927), .C(n1903), .Y(n6166) );
  NAND2X1 U3612 ( .A(ram[1729]), .B(n12927), .Y(n1903) );
  OAI21X1 U3613 ( .A(n12764), .B(n12927), .C(n1904), .Y(n6167) );
  NAND2X1 U3614 ( .A(ram[1730]), .B(n12927), .Y(n1904) );
  OAI21X1 U3615 ( .A(n12758), .B(n12927), .C(n1905), .Y(n6168) );
  NAND2X1 U3616 ( .A(ram[1731]), .B(n12927), .Y(n1905) );
  OAI21X1 U3617 ( .A(n12752), .B(n12927), .C(n1906), .Y(n6169) );
  NAND2X1 U3618 ( .A(ram[1732]), .B(n12927), .Y(n1906) );
  OAI21X1 U3619 ( .A(n12746), .B(n12927), .C(n1907), .Y(n6170) );
  NAND2X1 U3620 ( .A(ram[1733]), .B(n12927), .Y(n1907) );
  OAI21X1 U3621 ( .A(n12740), .B(n12927), .C(n1908), .Y(n6171) );
  NAND2X1 U3622 ( .A(ram[1734]), .B(n12927), .Y(n1908) );
  OAI21X1 U3623 ( .A(n12734), .B(n12927), .C(n1909), .Y(n6172) );
  NAND2X1 U3624 ( .A(ram[1735]), .B(n12927), .Y(n1909) );
  OAI21X1 U3625 ( .A(n12728), .B(n12927), .C(n1910), .Y(n6173) );
  NAND2X1 U3626 ( .A(ram[1736]), .B(n12927), .Y(n1910) );
  OAI21X1 U3627 ( .A(n12722), .B(n12927), .C(n1911), .Y(n6174) );
  NAND2X1 U3628 ( .A(ram[1737]), .B(n12927), .Y(n1911) );
  OAI21X1 U3629 ( .A(n12716), .B(n12927), .C(n1912), .Y(n6175) );
  NAND2X1 U3630 ( .A(ram[1738]), .B(n12927), .Y(n1912) );
  OAI21X1 U3631 ( .A(n12710), .B(n12927), .C(n1913), .Y(n6176) );
  NAND2X1 U3632 ( .A(ram[1739]), .B(n12927), .Y(n1913) );
  OAI21X1 U3633 ( .A(n12704), .B(n12927), .C(n1914), .Y(n6177) );
  NAND2X1 U3634 ( .A(ram[1740]), .B(n12927), .Y(n1914) );
  OAI21X1 U3635 ( .A(n12698), .B(n12927), .C(n1915), .Y(n6178) );
  NAND2X1 U3636 ( .A(ram[1741]), .B(n12927), .Y(n1915) );
  OAI21X1 U3637 ( .A(n12694), .B(n12927), .C(n1916), .Y(n6179) );
  NAND2X1 U3638 ( .A(ram[1742]), .B(n12927), .Y(n1916) );
  OAI21X1 U3639 ( .A(n12688), .B(n12927), .C(n1917), .Y(n6180) );
  NAND2X1 U3640 ( .A(ram[1743]), .B(n12927), .Y(n1917) );
  OAI21X1 U3642 ( .A(n12777), .B(n12926), .C(n1919), .Y(n6181) );
  NAND2X1 U3643 ( .A(ram[1744]), .B(n12926), .Y(n1919) );
  OAI21X1 U3644 ( .A(n12771), .B(n12926), .C(n1920), .Y(n6182) );
  NAND2X1 U3645 ( .A(ram[1745]), .B(n12926), .Y(n1920) );
  OAI21X1 U3646 ( .A(n12763), .B(n12926), .C(n1921), .Y(n6183) );
  NAND2X1 U3647 ( .A(ram[1746]), .B(n12926), .Y(n1921) );
  OAI21X1 U3648 ( .A(n12757), .B(n12926), .C(n1922), .Y(n6184) );
  NAND2X1 U3649 ( .A(ram[1747]), .B(n12926), .Y(n1922) );
  OAI21X1 U3650 ( .A(n12751), .B(n12926), .C(n1923), .Y(n6185) );
  NAND2X1 U3651 ( .A(ram[1748]), .B(n12926), .Y(n1923) );
  OAI21X1 U3652 ( .A(n12745), .B(n12926), .C(n1924), .Y(n6186) );
  NAND2X1 U3653 ( .A(ram[1749]), .B(n12926), .Y(n1924) );
  OAI21X1 U3654 ( .A(n12739), .B(n12926), .C(n1925), .Y(n6187) );
  NAND2X1 U3655 ( .A(ram[1750]), .B(n12926), .Y(n1925) );
  OAI21X1 U3656 ( .A(n12733), .B(n12926), .C(n1926), .Y(n6188) );
  NAND2X1 U3657 ( .A(ram[1751]), .B(n12926), .Y(n1926) );
  OAI21X1 U3658 ( .A(n12727), .B(n12926), .C(n1927), .Y(n6189) );
  NAND2X1 U3659 ( .A(ram[1752]), .B(n12926), .Y(n1927) );
  OAI21X1 U3660 ( .A(n12721), .B(n12926), .C(n1928), .Y(n6190) );
  NAND2X1 U3661 ( .A(ram[1753]), .B(n12926), .Y(n1928) );
  OAI21X1 U3662 ( .A(n12715), .B(n12926), .C(n1929), .Y(n6191) );
  NAND2X1 U3663 ( .A(ram[1754]), .B(n12926), .Y(n1929) );
  OAI21X1 U3664 ( .A(n12709), .B(n12926), .C(n1930), .Y(n6192) );
  NAND2X1 U3665 ( .A(ram[1755]), .B(n12926), .Y(n1930) );
  OAI21X1 U3666 ( .A(n12703), .B(n12926), .C(n1931), .Y(n6193) );
  NAND2X1 U3667 ( .A(ram[1756]), .B(n12926), .Y(n1931) );
  OAI21X1 U3668 ( .A(n12697), .B(n12926), .C(n1932), .Y(n6194) );
  NAND2X1 U3669 ( .A(ram[1757]), .B(n12926), .Y(n1932) );
  OAI21X1 U3670 ( .A(n12693), .B(n12926), .C(n1933), .Y(n6195) );
  NAND2X1 U3671 ( .A(ram[1758]), .B(n12926), .Y(n1933) );
  OAI21X1 U3672 ( .A(n12687), .B(n12926), .C(n1934), .Y(n6196) );
  NAND2X1 U3673 ( .A(ram[1759]), .B(n12926), .Y(n1934) );
  OAI21X1 U3675 ( .A(n13071), .B(n12925), .C(n1936), .Y(n6197) );
  NAND2X1 U3676 ( .A(ram[1760]), .B(n12925), .Y(n1936) );
  OAI21X1 U3677 ( .A(n13070), .B(n12925), .C(n1937), .Y(n6198) );
  NAND2X1 U3678 ( .A(ram[1761]), .B(n12925), .Y(n1937) );
  OAI21X1 U3679 ( .A(n12765), .B(n12925), .C(n1938), .Y(n6199) );
  NAND2X1 U3680 ( .A(ram[1762]), .B(n12925), .Y(n1938) );
  OAI21X1 U3681 ( .A(n12759), .B(n12925), .C(n1939), .Y(n6200) );
  NAND2X1 U3682 ( .A(ram[1763]), .B(n12925), .Y(n1939) );
  OAI21X1 U3683 ( .A(n12753), .B(n12925), .C(n1940), .Y(n6201) );
  NAND2X1 U3684 ( .A(ram[1764]), .B(n12925), .Y(n1940) );
  OAI21X1 U3685 ( .A(n12747), .B(n12925), .C(n1941), .Y(n6202) );
  NAND2X1 U3686 ( .A(ram[1765]), .B(n12925), .Y(n1941) );
  OAI21X1 U3687 ( .A(n12741), .B(n12925), .C(n1942), .Y(n6203) );
  NAND2X1 U3688 ( .A(ram[1766]), .B(n12925), .Y(n1942) );
  OAI21X1 U3689 ( .A(n12735), .B(n12925), .C(n1943), .Y(n6204) );
  NAND2X1 U3690 ( .A(ram[1767]), .B(n12925), .Y(n1943) );
  OAI21X1 U3691 ( .A(n12729), .B(n12925), .C(n1944), .Y(n6205) );
  NAND2X1 U3692 ( .A(ram[1768]), .B(n12925), .Y(n1944) );
  OAI21X1 U3693 ( .A(n12723), .B(n12925), .C(n1945), .Y(n6206) );
  NAND2X1 U3694 ( .A(ram[1769]), .B(n12925), .Y(n1945) );
  OAI21X1 U3695 ( .A(n12717), .B(n12925), .C(n1946), .Y(n6207) );
  NAND2X1 U3696 ( .A(ram[1770]), .B(n12925), .Y(n1946) );
  OAI21X1 U3697 ( .A(n12711), .B(n12925), .C(n1947), .Y(n6208) );
  NAND2X1 U3698 ( .A(ram[1771]), .B(n12925), .Y(n1947) );
  OAI21X1 U3699 ( .A(n12705), .B(n12925), .C(n1948), .Y(n6209) );
  NAND2X1 U3700 ( .A(ram[1772]), .B(n12925), .Y(n1948) );
  OAI21X1 U3701 ( .A(n12699), .B(n12925), .C(n1949), .Y(n6210) );
  NAND2X1 U3702 ( .A(ram[1773]), .B(n12925), .Y(n1949) );
  OAI21X1 U3703 ( .A(n13057), .B(n12925), .C(n1950), .Y(n6211) );
  NAND2X1 U3704 ( .A(ram[1774]), .B(n12925), .Y(n1950) );
  OAI21X1 U3705 ( .A(n13056), .B(n12925), .C(n1951), .Y(n6212) );
  NAND2X1 U3706 ( .A(ram[1775]), .B(n12925), .Y(n1951) );
  OAI21X1 U3708 ( .A(n12775), .B(n12924), .C(n1953), .Y(n6213) );
  NAND2X1 U3709 ( .A(ram[1776]), .B(n12924), .Y(n1953) );
  OAI21X1 U3710 ( .A(n12769), .B(n12924), .C(n1954), .Y(n6214) );
  NAND2X1 U3711 ( .A(ram[1777]), .B(n12924), .Y(n1954) );
  OAI21X1 U3712 ( .A(n12765), .B(n12924), .C(n1955), .Y(n6215) );
  NAND2X1 U3713 ( .A(ram[1778]), .B(n12924), .Y(n1955) );
  OAI21X1 U3714 ( .A(n12759), .B(n12924), .C(n1956), .Y(n6216) );
  NAND2X1 U3715 ( .A(ram[1779]), .B(n12924), .Y(n1956) );
  OAI21X1 U3716 ( .A(n12753), .B(n12924), .C(n1957), .Y(n6217) );
  NAND2X1 U3717 ( .A(ram[1780]), .B(n12924), .Y(n1957) );
  OAI21X1 U3718 ( .A(n12747), .B(n12924), .C(n1958), .Y(n6218) );
  NAND2X1 U3719 ( .A(ram[1781]), .B(n12924), .Y(n1958) );
  OAI21X1 U3720 ( .A(n12741), .B(n12924), .C(n1959), .Y(n6219) );
  NAND2X1 U3721 ( .A(ram[1782]), .B(n12924), .Y(n1959) );
  OAI21X1 U3722 ( .A(n12735), .B(n12924), .C(n1960), .Y(n6220) );
  NAND2X1 U3723 ( .A(ram[1783]), .B(n12924), .Y(n1960) );
  OAI21X1 U3724 ( .A(n12729), .B(n12924), .C(n1961), .Y(n6221) );
  NAND2X1 U3725 ( .A(ram[1784]), .B(n12924), .Y(n1961) );
  OAI21X1 U3726 ( .A(n12723), .B(n12924), .C(n1962), .Y(n6222) );
  NAND2X1 U3727 ( .A(ram[1785]), .B(n12924), .Y(n1962) );
  OAI21X1 U3728 ( .A(n12717), .B(n12924), .C(n1963), .Y(n6223) );
  NAND2X1 U3729 ( .A(ram[1786]), .B(n12924), .Y(n1963) );
  OAI21X1 U3730 ( .A(n12711), .B(n12924), .C(n1964), .Y(n6224) );
  NAND2X1 U3731 ( .A(ram[1787]), .B(n12924), .Y(n1964) );
  OAI21X1 U3732 ( .A(n12705), .B(n12924), .C(n1965), .Y(n6225) );
  NAND2X1 U3733 ( .A(ram[1788]), .B(n12924), .Y(n1965) );
  OAI21X1 U3734 ( .A(n12699), .B(n12924), .C(n1966), .Y(n6226) );
  NAND2X1 U3735 ( .A(ram[1789]), .B(n12924), .Y(n1966) );
  OAI21X1 U3736 ( .A(n12691), .B(n12924), .C(n1967), .Y(n6227) );
  NAND2X1 U3737 ( .A(ram[1790]), .B(n12924), .Y(n1967) );
  OAI21X1 U3738 ( .A(n12685), .B(n12924), .C(n1968), .Y(n6228) );
  NAND2X1 U3739 ( .A(ram[1791]), .B(n12924), .Y(n1968) );
  NAND3X1 U3741 ( .A(n875), .B(mem_write_en), .C(n1423), .Y(n1969) );
  OAI21X1 U3742 ( .A(n12779), .B(n12923), .C(n1971), .Y(n6229) );
  NAND2X1 U3743 ( .A(ram[1792]), .B(n12923), .Y(n1971) );
  OAI21X1 U3744 ( .A(n12773), .B(n12923), .C(n1972), .Y(n6230) );
  NAND2X1 U3745 ( .A(ram[1793]), .B(n12923), .Y(n1972) );
  OAI21X1 U3746 ( .A(n12762), .B(n12923), .C(n1973), .Y(n6231) );
  NAND2X1 U3747 ( .A(ram[1794]), .B(n12923), .Y(n1973) );
  OAI21X1 U3748 ( .A(n12756), .B(n12923), .C(n1974), .Y(n6232) );
  NAND2X1 U3749 ( .A(ram[1795]), .B(n12923), .Y(n1974) );
  OAI21X1 U3750 ( .A(n12750), .B(n12923), .C(n1975), .Y(n6233) );
  NAND2X1 U3751 ( .A(ram[1796]), .B(n12923), .Y(n1975) );
  OAI21X1 U3752 ( .A(n12744), .B(n12923), .C(n1976), .Y(n6234) );
  NAND2X1 U3753 ( .A(ram[1797]), .B(n12923), .Y(n1976) );
  OAI21X1 U3754 ( .A(n12738), .B(n12923), .C(n1977), .Y(n6235) );
  NAND2X1 U3755 ( .A(ram[1798]), .B(n12923), .Y(n1977) );
  OAI21X1 U3756 ( .A(n12732), .B(n12923), .C(n1978), .Y(n6236) );
  NAND2X1 U3757 ( .A(ram[1799]), .B(n12923), .Y(n1978) );
  OAI21X1 U3758 ( .A(n12726), .B(n12923), .C(n1979), .Y(n6237) );
  NAND2X1 U3759 ( .A(ram[1800]), .B(n12923), .Y(n1979) );
  OAI21X1 U3760 ( .A(n12720), .B(n12923), .C(n1980), .Y(n6238) );
  NAND2X1 U3761 ( .A(ram[1801]), .B(n12923), .Y(n1980) );
  OAI21X1 U3762 ( .A(n12714), .B(n12923), .C(n1981), .Y(n6239) );
  NAND2X1 U3763 ( .A(ram[1802]), .B(n12923), .Y(n1981) );
  OAI21X1 U3764 ( .A(n12708), .B(n12923), .C(n1982), .Y(n6240) );
  NAND2X1 U3765 ( .A(ram[1803]), .B(n12923), .Y(n1982) );
  OAI21X1 U3766 ( .A(n12702), .B(n12923), .C(n1983), .Y(n6241) );
  NAND2X1 U3767 ( .A(ram[1804]), .B(n12923), .Y(n1983) );
  OAI21X1 U3768 ( .A(n12696), .B(n12923), .C(n1984), .Y(n6242) );
  NAND2X1 U3769 ( .A(ram[1805]), .B(n12923), .Y(n1984) );
  OAI21X1 U3770 ( .A(n12695), .B(n12923), .C(n1985), .Y(n6243) );
  NAND2X1 U3771 ( .A(ram[1806]), .B(n12923), .Y(n1985) );
  OAI21X1 U3772 ( .A(n12689), .B(n12923), .C(n1986), .Y(n6244) );
  NAND2X1 U3773 ( .A(ram[1807]), .B(n12923), .Y(n1986) );
  OAI21X1 U3775 ( .A(n12779), .B(n12922), .C(n1988), .Y(n6245) );
  NAND2X1 U3776 ( .A(ram[1808]), .B(n12922), .Y(n1988) );
  OAI21X1 U3777 ( .A(n12773), .B(n12922), .C(n1989), .Y(n6246) );
  NAND2X1 U3778 ( .A(ram[1809]), .B(n12922), .Y(n1989) );
  OAI21X1 U3779 ( .A(n12767), .B(n12922), .C(n1990), .Y(n6247) );
  NAND2X1 U3780 ( .A(ram[1810]), .B(n12922), .Y(n1990) );
  OAI21X1 U3781 ( .A(n12761), .B(n12922), .C(n1991), .Y(n6248) );
  NAND2X1 U3782 ( .A(ram[1811]), .B(n12922), .Y(n1991) );
  OAI21X1 U3783 ( .A(n12755), .B(n12922), .C(n1992), .Y(n6249) );
  NAND2X1 U3784 ( .A(ram[1812]), .B(n12922), .Y(n1992) );
  OAI21X1 U3785 ( .A(n12749), .B(n12922), .C(n1993), .Y(n6250) );
  NAND2X1 U3786 ( .A(ram[1813]), .B(n12922), .Y(n1993) );
  OAI21X1 U3787 ( .A(n12743), .B(n12922), .C(n1994), .Y(n6251) );
  NAND2X1 U3788 ( .A(ram[1814]), .B(n12922), .Y(n1994) );
  OAI21X1 U3789 ( .A(n12737), .B(n12922), .C(n1995), .Y(n6252) );
  NAND2X1 U3790 ( .A(ram[1815]), .B(n12922), .Y(n1995) );
  OAI21X1 U3791 ( .A(n12731), .B(n12922), .C(n1996), .Y(n6253) );
  NAND2X1 U3792 ( .A(ram[1816]), .B(n12922), .Y(n1996) );
  OAI21X1 U3793 ( .A(n12725), .B(n12922), .C(n1997), .Y(n6254) );
  NAND2X1 U3794 ( .A(ram[1817]), .B(n12922), .Y(n1997) );
  OAI21X1 U3795 ( .A(n12719), .B(n12922), .C(n1998), .Y(n6255) );
  NAND2X1 U3796 ( .A(ram[1818]), .B(n12922), .Y(n1998) );
  OAI21X1 U3797 ( .A(n12713), .B(n12922), .C(n1999), .Y(n6256) );
  NAND2X1 U3798 ( .A(ram[1819]), .B(n12922), .Y(n1999) );
  OAI21X1 U3799 ( .A(n12707), .B(n12922), .C(n2000), .Y(n6257) );
  NAND2X1 U3800 ( .A(ram[1820]), .B(n12922), .Y(n2000) );
  OAI21X1 U3801 ( .A(n12701), .B(n12922), .C(n2001), .Y(n6258) );
  NAND2X1 U3802 ( .A(ram[1821]), .B(n12922), .Y(n2001) );
  OAI21X1 U3803 ( .A(n12695), .B(n12922), .C(n2002), .Y(n6259) );
  NAND2X1 U3804 ( .A(ram[1822]), .B(n12922), .Y(n2002) );
  OAI21X1 U3805 ( .A(n12689), .B(n12922), .C(n2003), .Y(n6260) );
  NAND2X1 U3806 ( .A(ram[1823]), .B(n12922), .Y(n2003) );
  OAI21X1 U3808 ( .A(n12774), .B(n12921), .C(n2005), .Y(n6261) );
  NAND2X1 U3809 ( .A(ram[1824]), .B(n12921), .Y(n2005) );
  OAI21X1 U3810 ( .A(n12768), .B(n12921), .C(n2006), .Y(n6262) );
  NAND2X1 U3811 ( .A(ram[1825]), .B(n12921), .Y(n2006) );
  OAI21X1 U3812 ( .A(n12764), .B(n12921), .C(n2007), .Y(n6263) );
  NAND2X1 U3813 ( .A(ram[1826]), .B(n12921), .Y(n2007) );
  OAI21X1 U3814 ( .A(n12758), .B(n12921), .C(n2008), .Y(n6264) );
  NAND2X1 U3815 ( .A(ram[1827]), .B(n12921), .Y(n2008) );
  OAI21X1 U3816 ( .A(n12752), .B(n12921), .C(n2009), .Y(n6265) );
  NAND2X1 U3817 ( .A(ram[1828]), .B(n12921), .Y(n2009) );
  OAI21X1 U3818 ( .A(n12746), .B(n12921), .C(n2010), .Y(n6266) );
  NAND2X1 U3819 ( .A(ram[1829]), .B(n12921), .Y(n2010) );
  OAI21X1 U3820 ( .A(n12740), .B(n12921), .C(n2011), .Y(n6267) );
  NAND2X1 U3821 ( .A(ram[1830]), .B(n12921), .Y(n2011) );
  OAI21X1 U3822 ( .A(n12734), .B(n12921), .C(n2012), .Y(n6268) );
  NAND2X1 U3823 ( .A(ram[1831]), .B(n12921), .Y(n2012) );
  OAI21X1 U3824 ( .A(n12728), .B(n12921), .C(n2013), .Y(n6269) );
  NAND2X1 U3825 ( .A(ram[1832]), .B(n12921), .Y(n2013) );
  OAI21X1 U3826 ( .A(n12722), .B(n12921), .C(n2014), .Y(n6270) );
  NAND2X1 U3827 ( .A(ram[1833]), .B(n12921), .Y(n2014) );
  OAI21X1 U3828 ( .A(n12716), .B(n12921), .C(n2015), .Y(n6271) );
  NAND2X1 U3829 ( .A(ram[1834]), .B(n12921), .Y(n2015) );
  OAI21X1 U3830 ( .A(n12710), .B(n12921), .C(n2016), .Y(n6272) );
  NAND2X1 U3831 ( .A(ram[1835]), .B(n12921), .Y(n2016) );
  OAI21X1 U3832 ( .A(n12704), .B(n12921), .C(n2017), .Y(n6273) );
  NAND2X1 U3833 ( .A(ram[1836]), .B(n12921), .Y(n2017) );
  OAI21X1 U3834 ( .A(n12698), .B(n12921), .C(n2018), .Y(n6274) );
  NAND2X1 U3835 ( .A(ram[1837]), .B(n12921), .Y(n2018) );
  OAI21X1 U3836 ( .A(n12690), .B(n12921), .C(n2019), .Y(n6275) );
  NAND2X1 U3837 ( .A(ram[1838]), .B(n12921), .Y(n2019) );
  OAI21X1 U3838 ( .A(n12684), .B(n12921), .C(n2020), .Y(n6276) );
  NAND2X1 U3839 ( .A(ram[1839]), .B(n12921), .Y(n2020) );
  OAI21X1 U3841 ( .A(n12776), .B(n12920), .C(n2022), .Y(n6277) );
  NAND2X1 U3842 ( .A(ram[1840]), .B(n12920), .Y(n2022) );
  OAI21X1 U3843 ( .A(n12770), .B(n12920), .C(n2023), .Y(n6278) );
  NAND2X1 U3844 ( .A(ram[1841]), .B(n12920), .Y(n2023) );
  OAI21X1 U3845 ( .A(n12766), .B(n12920), .C(n2024), .Y(n6279) );
  NAND2X1 U3846 ( .A(ram[1842]), .B(n12920), .Y(n2024) );
  OAI21X1 U3847 ( .A(n12760), .B(n12920), .C(n2025), .Y(n6280) );
  NAND2X1 U3848 ( .A(ram[1843]), .B(n12920), .Y(n2025) );
  OAI21X1 U3849 ( .A(n12754), .B(n12920), .C(n2026), .Y(n6281) );
  NAND2X1 U3850 ( .A(ram[1844]), .B(n12920), .Y(n2026) );
  OAI21X1 U3851 ( .A(n12748), .B(n12920), .C(n2027), .Y(n6282) );
  NAND2X1 U3852 ( .A(ram[1845]), .B(n12920), .Y(n2027) );
  OAI21X1 U3853 ( .A(n12742), .B(n12920), .C(n2028), .Y(n6283) );
  NAND2X1 U3854 ( .A(ram[1846]), .B(n12920), .Y(n2028) );
  OAI21X1 U3855 ( .A(n12736), .B(n12920), .C(n2029), .Y(n6284) );
  NAND2X1 U3856 ( .A(ram[1847]), .B(n12920), .Y(n2029) );
  OAI21X1 U3857 ( .A(n12730), .B(n12920), .C(n2030), .Y(n6285) );
  NAND2X1 U3858 ( .A(ram[1848]), .B(n12920), .Y(n2030) );
  OAI21X1 U3859 ( .A(n12724), .B(n12920), .C(n2031), .Y(n6286) );
  NAND2X1 U3860 ( .A(ram[1849]), .B(n12920), .Y(n2031) );
  OAI21X1 U3861 ( .A(n12718), .B(n12920), .C(n2032), .Y(n6287) );
  NAND2X1 U3862 ( .A(ram[1850]), .B(n12920), .Y(n2032) );
  OAI21X1 U3863 ( .A(n12712), .B(n12920), .C(n2033), .Y(n6288) );
  NAND2X1 U3864 ( .A(ram[1851]), .B(n12920), .Y(n2033) );
  OAI21X1 U3865 ( .A(n12706), .B(n12920), .C(n2034), .Y(n6289) );
  NAND2X1 U3866 ( .A(ram[1852]), .B(n12920), .Y(n2034) );
  OAI21X1 U3867 ( .A(n12700), .B(n12920), .C(n2035), .Y(n6290) );
  NAND2X1 U3868 ( .A(ram[1853]), .B(n12920), .Y(n2035) );
  OAI21X1 U3869 ( .A(n12692), .B(n12920), .C(n2036), .Y(n6291) );
  NAND2X1 U3870 ( .A(ram[1854]), .B(n12920), .Y(n2036) );
  OAI21X1 U3871 ( .A(n12686), .B(n12920), .C(n2037), .Y(n6292) );
  NAND2X1 U3872 ( .A(ram[1855]), .B(n12920), .Y(n2037) );
  OAI21X1 U3874 ( .A(n12776), .B(n12919), .C(n2039), .Y(n6293) );
  NAND2X1 U3875 ( .A(ram[1856]), .B(n12919), .Y(n2039) );
  OAI21X1 U3876 ( .A(n12770), .B(n12919), .C(n2040), .Y(n6294) );
  NAND2X1 U3877 ( .A(ram[1857]), .B(n12919), .Y(n2040) );
  OAI21X1 U3878 ( .A(n12765), .B(n12919), .C(n2041), .Y(n6295) );
  NAND2X1 U3879 ( .A(ram[1858]), .B(n12919), .Y(n2041) );
  OAI21X1 U3880 ( .A(n12759), .B(n12919), .C(n2042), .Y(n6296) );
  NAND2X1 U3881 ( .A(ram[1859]), .B(n12919), .Y(n2042) );
  OAI21X1 U3882 ( .A(n12753), .B(n12919), .C(n2043), .Y(n6297) );
  NAND2X1 U3883 ( .A(ram[1860]), .B(n12919), .Y(n2043) );
  OAI21X1 U3884 ( .A(n12747), .B(n12919), .C(n2044), .Y(n6298) );
  NAND2X1 U3885 ( .A(ram[1861]), .B(n12919), .Y(n2044) );
  OAI21X1 U3886 ( .A(n12741), .B(n12919), .C(n2045), .Y(n6299) );
  NAND2X1 U3887 ( .A(ram[1862]), .B(n12919), .Y(n2045) );
  OAI21X1 U3888 ( .A(n12735), .B(n12919), .C(n2046), .Y(n6300) );
  NAND2X1 U3889 ( .A(ram[1863]), .B(n12919), .Y(n2046) );
  OAI21X1 U3890 ( .A(n12729), .B(n12919), .C(n2047), .Y(n6301) );
  NAND2X1 U3891 ( .A(ram[1864]), .B(n12919), .Y(n2047) );
  OAI21X1 U3892 ( .A(n12723), .B(n12919), .C(n2048), .Y(n6302) );
  NAND2X1 U3893 ( .A(ram[1865]), .B(n12919), .Y(n2048) );
  OAI21X1 U3894 ( .A(n12717), .B(n12919), .C(n2049), .Y(n6303) );
  NAND2X1 U3895 ( .A(ram[1866]), .B(n12919), .Y(n2049) );
  OAI21X1 U3896 ( .A(n12711), .B(n12919), .C(n2050), .Y(n6304) );
  NAND2X1 U3897 ( .A(ram[1867]), .B(n12919), .Y(n2050) );
  OAI21X1 U3898 ( .A(n12705), .B(n12919), .C(n2051), .Y(n6305) );
  NAND2X1 U3899 ( .A(ram[1868]), .B(n12919), .Y(n2051) );
  OAI21X1 U3900 ( .A(n12699), .B(n12919), .C(n2052), .Y(n6306) );
  NAND2X1 U3901 ( .A(ram[1869]), .B(n12919), .Y(n2052) );
  OAI21X1 U3902 ( .A(n12692), .B(n12919), .C(n2053), .Y(n6307) );
  NAND2X1 U3903 ( .A(ram[1870]), .B(n12919), .Y(n2053) );
  OAI21X1 U3904 ( .A(n12686), .B(n12919), .C(n2054), .Y(n6308) );
  NAND2X1 U3905 ( .A(ram[1871]), .B(n12919), .Y(n2054) );
  OAI21X1 U3907 ( .A(n12775), .B(n12918), .C(n2056), .Y(n6309) );
  NAND2X1 U3908 ( .A(ram[1872]), .B(n12918), .Y(n2056) );
  OAI21X1 U3909 ( .A(n12769), .B(n12918), .C(n2057), .Y(n6310) );
  NAND2X1 U3910 ( .A(ram[1873]), .B(n12918), .Y(n2057) );
  OAI21X1 U3911 ( .A(n12762), .B(n12918), .C(n2058), .Y(n6311) );
  NAND2X1 U3912 ( .A(ram[1874]), .B(n12918), .Y(n2058) );
  OAI21X1 U3913 ( .A(n12756), .B(n12918), .C(n2059), .Y(n6312) );
  NAND2X1 U3914 ( .A(ram[1875]), .B(n12918), .Y(n2059) );
  OAI21X1 U3915 ( .A(n12750), .B(n12918), .C(n2060), .Y(n6313) );
  NAND2X1 U3916 ( .A(ram[1876]), .B(n12918), .Y(n2060) );
  OAI21X1 U3917 ( .A(n12744), .B(n12918), .C(n2061), .Y(n6314) );
  NAND2X1 U3918 ( .A(ram[1877]), .B(n12918), .Y(n2061) );
  OAI21X1 U3919 ( .A(n12738), .B(n12918), .C(n2062), .Y(n6315) );
  NAND2X1 U3920 ( .A(ram[1878]), .B(n12918), .Y(n2062) );
  OAI21X1 U3921 ( .A(n12732), .B(n12918), .C(n2063), .Y(n6316) );
  NAND2X1 U3922 ( .A(ram[1879]), .B(n12918), .Y(n2063) );
  OAI21X1 U3923 ( .A(n12726), .B(n12918), .C(n2064), .Y(n6317) );
  NAND2X1 U3924 ( .A(ram[1880]), .B(n12918), .Y(n2064) );
  OAI21X1 U3925 ( .A(n12720), .B(n12918), .C(n2065), .Y(n6318) );
  NAND2X1 U3926 ( .A(ram[1881]), .B(n12918), .Y(n2065) );
  OAI21X1 U3927 ( .A(n12714), .B(n12918), .C(n2066), .Y(n6319) );
  NAND2X1 U3928 ( .A(ram[1882]), .B(n12918), .Y(n2066) );
  OAI21X1 U3929 ( .A(n12708), .B(n12918), .C(n2067), .Y(n6320) );
  NAND2X1 U3930 ( .A(ram[1883]), .B(n12918), .Y(n2067) );
  OAI21X1 U3931 ( .A(n12702), .B(n12918), .C(n2068), .Y(n6321) );
  NAND2X1 U3932 ( .A(ram[1884]), .B(n12918), .Y(n2068) );
  OAI21X1 U3933 ( .A(n12696), .B(n12918), .C(n2069), .Y(n6322) );
  NAND2X1 U3934 ( .A(ram[1885]), .B(n12918), .Y(n2069) );
  OAI21X1 U3935 ( .A(n12691), .B(n12918), .C(n2070), .Y(n6323) );
  NAND2X1 U3936 ( .A(ram[1886]), .B(n12918), .Y(n2070) );
  OAI21X1 U3937 ( .A(n12685), .B(n12918), .C(n2071), .Y(n6324) );
  NAND2X1 U3938 ( .A(ram[1887]), .B(n12918), .Y(n2071) );
  OAI21X1 U3940 ( .A(n12774), .B(n12917), .C(n2073), .Y(n6325) );
  NAND2X1 U3941 ( .A(ram[1888]), .B(n12917), .Y(n2073) );
  OAI21X1 U3942 ( .A(n12768), .B(n12917), .C(n2074), .Y(n6326) );
  NAND2X1 U3943 ( .A(ram[1889]), .B(n12917), .Y(n2074) );
  OAI21X1 U3944 ( .A(n12763), .B(n12917), .C(n2075), .Y(n6327) );
  NAND2X1 U3945 ( .A(ram[1890]), .B(n12917), .Y(n2075) );
  OAI21X1 U3946 ( .A(n12757), .B(n12917), .C(n2076), .Y(n6328) );
  NAND2X1 U3947 ( .A(ram[1891]), .B(n12917), .Y(n2076) );
  OAI21X1 U3948 ( .A(n12751), .B(n12917), .C(n2077), .Y(n6329) );
  NAND2X1 U3949 ( .A(ram[1892]), .B(n12917), .Y(n2077) );
  OAI21X1 U3950 ( .A(n12745), .B(n12917), .C(n2078), .Y(n6330) );
  NAND2X1 U3951 ( .A(ram[1893]), .B(n12917), .Y(n2078) );
  OAI21X1 U3952 ( .A(n12739), .B(n12917), .C(n2079), .Y(n6331) );
  NAND2X1 U3953 ( .A(ram[1894]), .B(n12917), .Y(n2079) );
  OAI21X1 U3954 ( .A(n12733), .B(n12917), .C(n2080), .Y(n6332) );
  NAND2X1 U3955 ( .A(ram[1895]), .B(n12917), .Y(n2080) );
  OAI21X1 U3956 ( .A(n12727), .B(n12917), .C(n2081), .Y(n6333) );
  NAND2X1 U3957 ( .A(ram[1896]), .B(n12917), .Y(n2081) );
  OAI21X1 U3958 ( .A(n12721), .B(n12917), .C(n2082), .Y(n6334) );
  NAND2X1 U3959 ( .A(ram[1897]), .B(n12917), .Y(n2082) );
  OAI21X1 U3960 ( .A(n12715), .B(n12917), .C(n2083), .Y(n6335) );
  NAND2X1 U3961 ( .A(ram[1898]), .B(n12917), .Y(n2083) );
  OAI21X1 U3962 ( .A(n12709), .B(n12917), .C(n2084), .Y(n6336) );
  NAND2X1 U3963 ( .A(ram[1899]), .B(n12917), .Y(n2084) );
  OAI21X1 U3964 ( .A(n12703), .B(n12917), .C(n2085), .Y(n6337) );
  NAND2X1 U3965 ( .A(ram[1900]), .B(n12917), .Y(n2085) );
  OAI21X1 U3966 ( .A(n12697), .B(n12917), .C(n2086), .Y(n6338) );
  NAND2X1 U3967 ( .A(ram[1901]), .B(n12917), .Y(n2086) );
  OAI21X1 U3968 ( .A(n12690), .B(n12917), .C(n2087), .Y(n6339) );
  NAND2X1 U3969 ( .A(ram[1902]), .B(n12917), .Y(n2087) );
  OAI21X1 U3970 ( .A(n12684), .B(n12917), .C(n2088), .Y(n6340) );
  NAND2X1 U3971 ( .A(ram[1903]), .B(n12917), .Y(n2088) );
  OAI21X1 U3973 ( .A(n12774), .B(n12916), .C(n2090), .Y(n6341) );
  NAND2X1 U3974 ( .A(ram[1904]), .B(n12916), .Y(n2090) );
  OAI21X1 U3975 ( .A(n12768), .B(n12916), .C(n2091), .Y(n6342) );
  NAND2X1 U3976 ( .A(ram[1905]), .B(n12916), .Y(n2091) );
  OAI21X1 U3977 ( .A(n12763), .B(n12916), .C(n2092), .Y(n6343) );
  NAND2X1 U3978 ( .A(ram[1906]), .B(n12916), .Y(n2092) );
  OAI21X1 U3979 ( .A(n12757), .B(n12916), .C(n2093), .Y(n6344) );
  NAND2X1 U3980 ( .A(ram[1907]), .B(n12916), .Y(n2093) );
  OAI21X1 U3981 ( .A(n12751), .B(n12916), .C(n2094), .Y(n6345) );
  NAND2X1 U3982 ( .A(ram[1908]), .B(n12916), .Y(n2094) );
  OAI21X1 U3983 ( .A(n12745), .B(n12916), .C(n2095), .Y(n6346) );
  NAND2X1 U3984 ( .A(ram[1909]), .B(n12916), .Y(n2095) );
  OAI21X1 U3985 ( .A(n12739), .B(n12916), .C(n2096), .Y(n6347) );
  NAND2X1 U3986 ( .A(ram[1910]), .B(n12916), .Y(n2096) );
  OAI21X1 U3987 ( .A(n12733), .B(n12916), .C(n2097), .Y(n6348) );
  NAND2X1 U3988 ( .A(ram[1911]), .B(n12916), .Y(n2097) );
  OAI21X1 U3989 ( .A(n12727), .B(n12916), .C(n2098), .Y(n6349) );
  NAND2X1 U3990 ( .A(ram[1912]), .B(n12916), .Y(n2098) );
  OAI21X1 U3991 ( .A(n12721), .B(n12916), .C(n2099), .Y(n6350) );
  NAND2X1 U3992 ( .A(ram[1913]), .B(n12916), .Y(n2099) );
  OAI21X1 U3993 ( .A(n12715), .B(n12916), .C(n2100), .Y(n6351) );
  NAND2X1 U3994 ( .A(ram[1914]), .B(n12916), .Y(n2100) );
  OAI21X1 U3995 ( .A(n12709), .B(n12916), .C(n2101), .Y(n6352) );
  NAND2X1 U3996 ( .A(ram[1915]), .B(n12916), .Y(n2101) );
  OAI21X1 U3997 ( .A(n12703), .B(n12916), .C(n2102), .Y(n6353) );
  NAND2X1 U3998 ( .A(ram[1916]), .B(n12916), .Y(n2102) );
  OAI21X1 U3999 ( .A(n12697), .B(n12916), .C(n2103), .Y(n6354) );
  NAND2X1 U4000 ( .A(ram[1917]), .B(n12916), .Y(n2103) );
  OAI21X1 U4001 ( .A(n12690), .B(n12916), .C(n2104), .Y(n6355) );
  NAND2X1 U4002 ( .A(ram[1918]), .B(n12916), .Y(n2104) );
  OAI21X1 U4003 ( .A(n12684), .B(n12916), .C(n2105), .Y(n6356) );
  NAND2X1 U4004 ( .A(ram[1919]), .B(n12916), .Y(n2105) );
  OAI21X1 U4006 ( .A(n12776), .B(n12915), .C(n2107), .Y(n6357) );
  NAND2X1 U4007 ( .A(ram[1920]), .B(n12915), .Y(n2107) );
  OAI21X1 U4008 ( .A(n12770), .B(n12915), .C(n2108), .Y(n6358) );
  NAND2X1 U4009 ( .A(ram[1921]), .B(n12915), .Y(n2108) );
  OAI21X1 U4010 ( .A(n12762), .B(n12915), .C(n2109), .Y(n6359) );
  NAND2X1 U4011 ( .A(ram[1922]), .B(n12915), .Y(n2109) );
  OAI21X1 U4012 ( .A(n12756), .B(n12915), .C(n2110), .Y(n6360) );
  NAND2X1 U4013 ( .A(ram[1923]), .B(n12915), .Y(n2110) );
  OAI21X1 U4014 ( .A(n12750), .B(n12915), .C(n2111), .Y(n6361) );
  NAND2X1 U4015 ( .A(ram[1924]), .B(n12915), .Y(n2111) );
  OAI21X1 U4016 ( .A(n12744), .B(n12915), .C(n2112), .Y(n6362) );
  NAND2X1 U4017 ( .A(ram[1925]), .B(n12915), .Y(n2112) );
  OAI21X1 U4018 ( .A(n12738), .B(n12915), .C(n2113), .Y(n6363) );
  NAND2X1 U4019 ( .A(ram[1926]), .B(n12915), .Y(n2113) );
  OAI21X1 U4020 ( .A(n12732), .B(n12915), .C(n2114), .Y(n6364) );
  NAND2X1 U4021 ( .A(ram[1927]), .B(n12915), .Y(n2114) );
  OAI21X1 U4022 ( .A(n12726), .B(n12915), .C(n2115), .Y(n6365) );
  NAND2X1 U4023 ( .A(ram[1928]), .B(n12915), .Y(n2115) );
  OAI21X1 U4024 ( .A(n12720), .B(n12915), .C(n2116), .Y(n6366) );
  NAND2X1 U4025 ( .A(ram[1929]), .B(n12915), .Y(n2116) );
  OAI21X1 U4026 ( .A(n12714), .B(n12915), .C(n2117), .Y(n6367) );
  NAND2X1 U4027 ( .A(ram[1930]), .B(n12915), .Y(n2117) );
  OAI21X1 U4028 ( .A(n12708), .B(n12915), .C(n2118), .Y(n6368) );
  NAND2X1 U4029 ( .A(ram[1931]), .B(n12915), .Y(n2118) );
  OAI21X1 U4030 ( .A(n12702), .B(n12915), .C(n2119), .Y(n6369) );
  NAND2X1 U4031 ( .A(ram[1932]), .B(n12915), .Y(n2119) );
  OAI21X1 U4032 ( .A(n12696), .B(n12915), .C(n2120), .Y(n6370) );
  NAND2X1 U4033 ( .A(ram[1933]), .B(n12915), .Y(n2120) );
  OAI21X1 U4034 ( .A(n12692), .B(n12915), .C(n2121), .Y(n6371) );
  NAND2X1 U4035 ( .A(ram[1934]), .B(n12915), .Y(n2121) );
  OAI21X1 U4036 ( .A(n12686), .B(n12915), .C(n2122), .Y(n6372) );
  NAND2X1 U4037 ( .A(ram[1935]), .B(n12915), .Y(n2122) );
  OAI21X1 U4039 ( .A(n12774), .B(n12914), .C(n2124), .Y(n6373) );
  NAND2X1 U4040 ( .A(ram[1936]), .B(n12914), .Y(n2124) );
  OAI21X1 U4041 ( .A(n12768), .B(n12914), .C(n2125), .Y(n6374) );
  NAND2X1 U4042 ( .A(ram[1937]), .B(n12914), .Y(n2125) );
  OAI21X1 U4043 ( .A(n12762), .B(n12914), .C(n2126), .Y(n6375) );
  NAND2X1 U4044 ( .A(ram[1938]), .B(n12914), .Y(n2126) );
  OAI21X1 U4045 ( .A(n12756), .B(n12914), .C(n2127), .Y(n6376) );
  NAND2X1 U4046 ( .A(ram[1939]), .B(n12914), .Y(n2127) );
  OAI21X1 U4047 ( .A(n12750), .B(n12914), .C(n2128), .Y(n6377) );
  NAND2X1 U4048 ( .A(ram[1940]), .B(n12914), .Y(n2128) );
  OAI21X1 U4049 ( .A(n12744), .B(n12914), .C(n2129), .Y(n6378) );
  NAND2X1 U4050 ( .A(ram[1941]), .B(n12914), .Y(n2129) );
  OAI21X1 U4051 ( .A(n12738), .B(n12914), .C(n2130), .Y(n6379) );
  NAND2X1 U4052 ( .A(ram[1942]), .B(n12914), .Y(n2130) );
  OAI21X1 U4053 ( .A(n12732), .B(n12914), .C(n2131), .Y(n6380) );
  NAND2X1 U4054 ( .A(ram[1943]), .B(n12914), .Y(n2131) );
  OAI21X1 U4055 ( .A(n12726), .B(n12914), .C(n2132), .Y(n6381) );
  NAND2X1 U4056 ( .A(ram[1944]), .B(n12914), .Y(n2132) );
  OAI21X1 U4057 ( .A(n12720), .B(n12914), .C(n2133), .Y(n6382) );
  NAND2X1 U4058 ( .A(ram[1945]), .B(n12914), .Y(n2133) );
  OAI21X1 U4059 ( .A(n12714), .B(n12914), .C(n2134), .Y(n6383) );
  NAND2X1 U4060 ( .A(ram[1946]), .B(n12914), .Y(n2134) );
  OAI21X1 U4061 ( .A(n12708), .B(n12914), .C(n2135), .Y(n6384) );
  NAND2X1 U4062 ( .A(ram[1947]), .B(n12914), .Y(n2135) );
  OAI21X1 U4063 ( .A(n12702), .B(n12914), .C(n2136), .Y(n6385) );
  NAND2X1 U4064 ( .A(ram[1948]), .B(n12914), .Y(n2136) );
  OAI21X1 U4065 ( .A(n12696), .B(n12914), .C(n2137), .Y(n6386) );
  NAND2X1 U4066 ( .A(ram[1949]), .B(n12914), .Y(n2137) );
  OAI21X1 U4067 ( .A(n12690), .B(n12914), .C(n2138), .Y(n6387) );
  NAND2X1 U4068 ( .A(ram[1950]), .B(n12914), .Y(n2138) );
  OAI21X1 U4069 ( .A(n12684), .B(n12914), .C(n2139), .Y(n6388) );
  NAND2X1 U4070 ( .A(ram[1951]), .B(n12914), .Y(n2139) );
  OAI21X1 U4072 ( .A(n12775), .B(n12913), .C(n2141), .Y(n6389) );
  NAND2X1 U4073 ( .A(ram[1952]), .B(n12913), .Y(n2141) );
  OAI21X1 U4074 ( .A(n12769), .B(n12913), .C(n2142), .Y(n6390) );
  NAND2X1 U4075 ( .A(ram[1953]), .B(n12913), .Y(n2142) );
  OAI21X1 U4076 ( .A(n12763), .B(n12913), .C(n2143), .Y(n6391) );
  NAND2X1 U4077 ( .A(ram[1954]), .B(n12913), .Y(n2143) );
  OAI21X1 U4078 ( .A(n12757), .B(n12913), .C(n2144), .Y(n6392) );
  NAND2X1 U4079 ( .A(ram[1955]), .B(n12913), .Y(n2144) );
  OAI21X1 U4080 ( .A(n12751), .B(n12913), .C(n2145), .Y(n6393) );
  NAND2X1 U4081 ( .A(ram[1956]), .B(n12913), .Y(n2145) );
  OAI21X1 U4082 ( .A(n12745), .B(n12913), .C(n2146), .Y(n6394) );
  NAND2X1 U4083 ( .A(ram[1957]), .B(n12913), .Y(n2146) );
  OAI21X1 U4084 ( .A(n12739), .B(n12913), .C(n2147), .Y(n6395) );
  NAND2X1 U4085 ( .A(ram[1958]), .B(n12913), .Y(n2147) );
  OAI21X1 U4086 ( .A(n12733), .B(n12913), .C(n2148), .Y(n6396) );
  NAND2X1 U4087 ( .A(ram[1959]), .B(n12913), .Y(n2148) );
  OAI21X1 U4088 ( .A(n12727), .B(n12913), .C(n2149), .Y(n6397) );
  NAND2X1 U4089 ( .A(ram[1960]), .B(n12913), .Y(n2149) );
  OAI21X1 U4090 ( .A(n12721), .B(n12913), .C(n2150), .Y(n6398) );
  NAND2X1 U4091 ( .A(ram[1961]), .B(n12913), .Y(n2150) );
  OAI21X1 U4092 ( .A(n12715), .B(n12913), .C(n2151), .Y(n6399) );
  NAND2X1 U4093 ( .A(ram[1962]), .B(n12913), .Y(n2151) );
  OAI21X1 U4094 ( .A(n12709), .B(n12913), .C(n2152), .Y(n6400) );
  NAND2X1 U4095 ( .A(ram[1963]), .B(n12913), .Y(n2152) );
  OAI21X1 U4096 ( .A(n12703), .B(n12913), .C(n2153), .Y(n6401) );
  NAND2X1 U4097 ( .A(ram[1964]), .B(n12913), .Y(n2153) );
  OAI21X1 U4098 ( .A(n12697), .B(n12913), .C(n2154), .Y(n6402) );
  NAND2X1 U4099 ( .A(ram[1965]), .B(n12913), .Y(n2154) );
  OAI21X1 U4100 ( .A(n12691), .B(n12913), .C(n2155), .Y(n6403) );
  NAND2X1 U4101 ( .A(ram[1966]), .B(n12913), .Y(n2155) );
  OAI21X1 U4102 ( .A(n12685), .B(n12913), .C(n2156), .Y(n6404) );
  NAND2X1 U4103 ( .A(ram[1967]), .B(n12913), .Y(n2156) );
  OAI21X1 U4105 ( .A(n12774), .B(n12912), .C(n2158), .Y(n6405) );
  NAND2X1 U4106 ( .A(ram[1968]), .B(n12912), .Y(n2158) );
  OAI21X1 U4107 ( .A(n12768), .B(n12912), .C(n2159), .Y(n6406) );
  NAND2X1 U4108 ( .A(ram[1969]), .B(n12912), .Y(n2159) );
  OAI21X1 U4109 ( .A(n12767), .B(n12912), .C(n2160), .Y(n6407) );
  NAND2X1 U4110 ( .A(ram[1970]), .B(n12912), .Y(n2160) );
  OAI21X1 U4111 ( .A(n12761), .B(n12912), .C(n2161), .Y(n6408) );
  NAND2X1 U4112 ( .A(ram[1971]), .B(n12912), .Y(n2161) );
  OAI21X1 U4113 ( .A(n12755), .B(n12912), .C(n2162), .Y(n6409) );
  NAND2X1 U4114 ( .A(ram[1972]), .B(n12912), .Y(n2162) );
  OAI21X1 U4115 ( .A(n12749), .B(n12912), .C(n2163), .Y(n6410) );
  NAND2X1 U4116 ( .A(ram[1973]), .B(n12912), .Y(n2163) );
  OAI21X1 U4117 ( .A(n12743), .B(n12912), .C(n2164), .Y(n6411) );
  NAND2X1 U4118 ( .A(ram[1974]), .B(n12912), .Y(n2164) );
  OAI21X1 U4119 ( .A(n12737), .B(n12912), .C(n2165), .Y(n6412) );
  NAND2X1 U4120 ( .A(ram[1975]), .B(n12912), .Y(n2165) );
  OAI21X1 U4121 ( .A(n12731), .B(n12912), .C(n2166), .Y(n6413) );
  NAND2X1 U4122 ( .A(ram[1976]), .B(n12912), .Y(n2166) );
  OAI21X1 U4123 ( .A(n12725), .B(n12912), .C(n2167), .Y(n6414) );
  NAND2X1 U4124 ( .A(ram[1977]), .B(n12912), .Y(n2167) );
  OAI21X1 U4125 ( .A(n12719), .B(n12912), .C(n2168), .Y(n6415) );
  NAND2X1 U4126 ( .A(ram[1978]), .B(n12912), .Y(n2168) );
  OAI21X1 U4127 ( .A(n12713), .B(n12912), .C(n2169), .Y(n6416) );
  NAND2X1 U4128 ( .A(ram[1979]), .B(n12912), .Y(n2169) );
  OAI21X1 U4129 ( .A(n12707), .B(n12912), .C(n2170), .Y(n6417) );
  NAND2X1 U4130 ( .A(ram[1980]), .B(n12912), .Y(n2170) );
  OAI21X1 U4131 ( .A(n12701), .B(n12912), .C(n2171), .Y(n6418) );
  NAND2X1 U4132 ( .A(ram[1981]), .B(n12912), .Y(n2171) );
  OAI21X1 U4133 ( .A(n12690), .B(n12912), .C(n2172), .Y(n6419) );
  NAND2X1 U4134 ( .A(ram[1982]), .B(n12912), .Y(n2172) );
  OAI21X1 U4135 ( .A(n12684), .B(n12912), .C(n2173), .Y(n6420) );
  NAND2X1 U4136 ( .A(ram[1983]), .B(n12912), .Y(n2173) );
  OAI21X1 U4138 ( .A(n12777), .B(n12911), .C(n2175), .Y(n6421) );
  NAND2X1 U4139 ( .A(ram[1984]), .B(n12911), .Y(n2175) );
  OAI21X1 U4140 ( .A(n12771), .B(n12911), .C(n2176), .Y(n6422) );
  NAND2X1 U4141 ( .A(ram[1985]), .B(n12911), .Y(n2176) );
  OAI21X1 U4142 ( .A(n12767), .B(n12911), .C(n2177), .Y(n6423) );
  NAND2X1 U4143 ( .A(ram[1986]), .B(n12911), .Y(n2177) );
  OAI21X1 U4144 ( .A(n12761), .B(n12911), .C(n2178), .Y(n6424) );
  NAND2X1 U4145 ( .A(ram[1987]), .B(n12911), .Y(n2178) );
  OAI21X1 U4146 ( .A(n12755), .B(n12911), .C(n2179), .Y(n6425) );
  NAND2X1 U4147 ( .A(ram[1988]), .B(n12911), .Y(n2179) );
  OAI21X1 U4148 ( .A(n12749), .B(n12911), .C(n2180), .Y(n6426) );
  NAND2X1 U4149 ( .A(ram[1989]), .B(n12911), .Y(n2180) );
  OAI21X1 U4150 ( .A(n12743), .B(n12911), .C(n2181), .Y(n6427) );
  NAND2X1 U4151 ( .A(ram[1990]), .B(n12911), .Y(n2181) );
  OAI21X1 U4152 ( .A(n12737), .B(n12911), .C(n2182), .Y(n6428) );
  NAND2X1 U4153 ( .A(ram[1991]), .B(n12911), .Y(n2182) );
  OAI21X1 U4154 ( .A(n12731), .B(n12911), .C(n2183), .Y(n6429) );
  NAND2X1 U4155 ( .A(ram[1992]), .B(n12911), .Y(n2183) );
  OAI21X1 U4156 ( .A(n12725), .B(n12911), .C(n2184), .Y(n6430) );
  NAND2X1 U4157 ( .A(ram[1993]), .B(n12911), .Y(n2184) );
  OAI21X1 U4158 ( .A(n12719), .B(n12911), .C(n2185), .Y(n6431) );
  NAND2X1 U4159 ( .A(ram[1994]), .B(n12911), .Y(n2185) );
  OAI21X1 U4160 ( .A(n12713), .B(n12911), .C(n2186), .Y(n6432) );
  NAND2X1 U4161 ( .A(ram[1995]), .B(n12911), .Y(n2186) );
  OAI21X1 U4162 ( .A(n12707), .B(n12911), .C(n2187), .Y(n6433) );
  NAND2X1 U4163 ( .A(ram[1996]), .B(n12911), .Y(n2187) );
  OAI21X1 U4164 ( .A(n12701), .B(n12911), .C(n2188), .Y(n6434) );
  NAND2X1 U4165 ( .A(ram[1997]), .B(n12911), .Y(n2188) );
  OAI21X1 U4166 ( .A(n12693), .B(n12911), .C(n2189), .Y(n6435) );
  NAND2X1 U4167 ( .A(ram[1998]), .B(n12911), .Y(n2189) );
  OAI21X1 U4168 ( .A(n12687), .B(n12911), .C(n2190), .Y(n6436) );
  NAND2X1 U4169 ( .A(ram[1999]), .B(n12911), .Y(n2190) );
  OAI21X1 U4171 ( .A(n12778), .B(n12910), .C(n2192), .Y(n6437) );
  NAND2X1 U4172 ( .A(ram[2000]), .B(n12910), .Y(n2192) );
  OAI21X1 U4173 ( .A(n12772), .B(n12910), .C(n2193), .Y(n6438) );
  NAND2X1 U4174 ( .A(ram[2001]), .B(n12910), .Y(n2193) );
  OAI21X1 U4175 ( .A(n12766), .B(n12910), .C(n2194), .Y(n6439) );
  NAND2X1 U4176 ( .A(ram[2002]), .B(n12910), .Y(n2194) );
  OAI21X1 U4177 ( .A(n12760), .B(n12910), .C(n2195), .Y(n6440) );
  NAND2X1 U4178 ( .A(ram[2003]), .B(n12910), .Y(n2195) );
  OAI21X1 U4179 ( .A(n12754), .B(n12910), .C(n2196), .Y(n6441) );
  NAND2X1 U4180 ( .A(ram[2004]), .B(n12910), .Y(n2196) );
  OAI21X1 U4181 ( .A(n12748), .B(n12910), .C(n2197), .Y(n6442) );
  NAND2X1 U4182 ( .A(ram[2005]), .B(n12910), .Y(n2197) );
  OAI21X1 U4183 ( .A(n12742), .B(n12910), .C(n2198), .Y(n6443) );
  NAND2X1 U4184 ( .A(ram[2006]), .B(n12910), .Y(n2198) );
  OAI21X1 U4185 ( .A(n12736), .B(n12910), .C(n2199), .Y(n6444) );
  NAND2X1 U4186 ( .A(ram[2007]), .B(n12910), .Y(n2199) );
  OAI21X1 U4187 ( .A(n12730), .B(n12910), .C(n2200), .Y(n6445) );
  NAND2X1 U4188 ( .A(ram[2008]), .B(n12910), .Y(n2200) );
  OAI21X1 U4189 ( .A(n12724), .B(n12910), .C(n2201), .Y(n6446) );
  NAND2X1 U4190 ( .A(ram[2009]), .B(n12910), .Y(n2201) );
  OAI21X1 U4191 ( .A(n12718), .B(n12910), .C(n2202), .Y(n6447) );
  NAND2X1 U4192 ( .A(ram[2010]), .B(n12910), .Y(n2202) );
  OAI21X1 U4193 ( .A(n12712), .B(n12910), .C(n2203), .Y(n6448) );
  NAND2X1 U4194 ( .A(ram[2011]), .B(n12910), .Y(n2203) );
  OAI21X1 U4195 ( .A(n12706), .B(n12910), .C(n2204), .Y(n6449) );
  NAND2X1 U4196 ( .A(ram[2012]), .B(n12910), .Y(n2204) );
  OAI21X1 U4197 ( .A(n12700), .B(n12910), .C(n2205), .Y(n6450) );
  NAND2X1 U4198 ( .A(ram[2013]), .B(n12910), .Y(n2205) );
  OAI21X1 U4199 ( .A(n12694), .B(n12910), .C(n2206), .Y(n6451) );
  NAND2X1 U4200 ( .A(ram[2014]), .B(n12910), .Y(n2206) );
  OAI21X1 U4201 ( .A(n12688), .B(n12910), .C(n2207), .Y(n6452) );
  NAND2X1 U4202 ( .A(ram[2015]), .B(n12910), .Y(n2207) );
  OAI21X1 U4204 ( .A(n12779), .B(n12909), .C(n2209), .Y(n6453) );
  NAND2X1 U4205 ( .A(ram[2016]), .B(n12909), .Y(n2209) );
  OAI21X1 U4206 ( .A(n12773), .B(n12909), .C(n2210), .Y(n6454) );
  NAND2X1 U4207 ( .A(ram[2017]), .B(n12909), .Y(n2210) );
  OAI21X1 U4208 ( .A(n12764), .B(n12909), .C(n2211), .Y(n6455) );
  NAND2X1 U4209 ( .A(ram[2018]), .B(n12909), .Y(n2211) );
  OAI21X1 U4210 ( .A(n12758), .B(n12909), .C(n2212), .Y(n6456) );
  NAND2X1 U4211 ( .A(ram[2019]), .B(n12909), .Y(n2212) );
  OAI21X1 U4212 ( .A(n12752), .B(n12909), .C(n2213), .Y(n6457) );
  NAND2X1 U4213 ( .A(ram[2020]), .B(n12909), .Y(n2213) );
  OAI21X1 U4214 ( .A(n12746), .B(n12909), .C(n2214), .Y(n6458) );
  NAND2X1 U4215 ( .A(ram[2021]), .B(n12909), .Y(n2214) );
  OAI21X1 U4216 ( .A(n12740), .B(n12909), .C(n2215), .Y(n6459) );
  NAND2X1 U4217 ( .A(ram[2022]), .B(n12909), .Y(n2215) );
  OAI21X1 U4218 ( .A(n12734), .B(n12909), .C(n2216), .Y(n6460) );
  NAND2X1 U4219 ( .A(ram[2023]), .B(n12909), .Y(n2216) );
  OAI21X1 U4220 ( .A(n12728), .B(n12909), .C(n2217), .Y(n6461) );
  NAND2X1 U4221 ( .A(ram[2024]), .B(n12909), .Y(n2217) );
  OAI21X1 U4222 ( .A(n12722), .B(n12909), .C(n2218), .Y(n6462) );
  NAND2X1 U4223 ( .A(ram[2025]), .B(n12909), .Y(n2218) );
  OAI21X1 U4224 ( .A(n12716), .B(n12909), .C(n2219), .Y(n6463) );
  NAND2X1 U4225 ( .A(ram[2026]), .B(n12909), .Y(n2219) );
  OAI21X1 U4226 ( .A(n12710), .B(n12909), .C(n2220), .Y(n6464) );
  NAND2X1 U4227 ( .A(ram[2027]), .B(n12909), .Y(n2220) );
  OAI21X1 U4228 ( .A(n12704), .B(n12909), .C(n2221), .Y(n6465) );
  NAND2X1 U4229 ( .A(ram[2028]), .B(n12909), .Y(n2221) );
  OAI21X1 U4230 ( .A(n12698), .B(n12909), .C(n2222), .Y(n6466) );
  NAND2X1 U4231 ( .A(ram[2029]), .B(n12909), .Y(n2222) );
  OAI21X1 U4232 ( .A(n12695), .B(n12909), .C(n2223), .Y(n6467) );
  NAND2X1 U4233 ( .A(ram[2030]), .B(n12909), .Y(n2223) );
  OAI21X1 U4234 ( .A(n12689), .B(n12909), .C(n2224), .Y(n6468) );
  NAND2X1 U4235 ( .A(ram[2031]), .B(n12909), .Y(n2224) );
  OAI21X1 U4237 ( .A(n12778), .B(n12908), .C(n2226), .Y(n6469) );
  NAND2X1 U4238 ( .A(ram[2032]), .B(n12908), .Y(n2226) );
  OAI21X1 U4239 ( .A(n12772), .B(n12908), .C(n2227), .Y(n6470) );
  NAND2X1 U4240 ( .A(ram[2033]), .B(n12908), .Y(n2227) );
  OAI21X1 U4241 ( .A(n12762), .B(n12908), .C(n2228), .Y(n6471) );
  NAND2X1 U4242 ( .A(ram[2034]), .B(n12908), .Y(n2228) );
  OAI21X1 U4243 ( .A(n12756), .B(n12908), .C(n2229), .Y(n6472) );
  NAND2X1 U4244 ( .A(ram[2035]), .B(n12908), .Y(n2229) );
  OAI21X1 U4245 ( .A(n12750), .B(n12908), .C(n2230), .Y(n6473) );
  NAND2X1 U4246 ( .A(ram[2036]), .B(n12908), .Y(n2230) );
  OAI21X1 U4247 ( .A(n12744), .B(n12908), .C(n2231), .Y(n6474) );
  NAND2X1 U4248 ( .A(ram[2037]), .B(n12908), .Y(n2231) );
  OAI21X1 U4249 ( .A(n12738), .B(n12908), .C(n2232), .Y(n6475) );
  NAND2X1 U4250 ( .A(ram[2038]), .B(n12908), .Y(n2232) );
  OAI21X1 U4251 ( .A(n12732), .B(n12908), .C(n2233), .Y(n6476) );
  NAND2X1 U4252 ( .A(ram[2039]), .B(n12908), .Y(n2233) );
  OAI21X1 U4253 ( .A(n12726), .B(n12908), .C(n2234), .Y(n6477) );
  NAND2X1 U4254 ( .A(ram[2040]), .B(n12908), .Y(n2234) );
  OAI21X1 U4255 ( .A(n12720), .B(n12908), .C(n2235), .Y(n6478) );
  NAND2X1 U4256 ( .A(ram[2041]), .B(n12908), .Y(n2235) );
  OAI21X1 U4257 ( .A(n12714), .B(n12908), .C(n2236), .Y(n6479) );
  NAND2X1 U4258 ( .A(ram[2042]), .B(n12908), .Y(n2236) );
  OAI21X1 U4259 ( .A(n12708), .B(n12908), .C(n2237), .Y(n6480) );
  NAND2X1 U4260 ( .A(ram[2043]), .B(n12908), .Y(n2237) );
  OAI21X1 U4261 ( .A(n12702), .B(n12908), .C(n2238), .Y(n6481) );
  NAND2X1 U4262 ( .A(ram[2044]), .B(n12908), .Y(n2238) );
  OAI21X1 U4263 ( .A(n12696), .B(n12908), .C(n2239), .Y(n6482) );
  NAND2X1 U4264 ( .A(ram[2045]), .B(n12908), .Y(n2239) );
  OAI21X1 U4265 ( .A(n12694), .B(n12908), .C(n2240), .Y(n6483) );
  NAND2X1 U4266 ( .A(ram[2046]), .B(n12908), .Y(n2240) );
  OAI21X1 U4267 ( .A(n12688), .B(n12908), .C(n2241), .Y(n6484) );
  NAND2X1 U4268 ( .A(ram[2047]), .B(n12908), .Y(n2241) );
  NAND3X1 U4270 ( .A(n1149), .B(mem_write_en), .C(n1423), .Y(n2242) );
  NOR2X1 U4271 ( .A(n13039), .B(mem_access_addr[7]), .Y(n1423) );
  OAI21X1 U4272 ( .A(n12777), .B(n12907), .C(n2244), .Y(n6485) );
  NAND2X1 U4273 ( .A(ram[2048]), .B(n12907), .Y(n2244) );
  OAI21X1 U4274 ( .A(n12771), .B(n12907), .C(n2245), .Y(n6486) );
  NAND2X1 U4275 ( .A(ram[2049]), .B(n12907), .Y(n2245) );
  OAI21X1 U4276 ( .A(n12767), .B(n12907), .C(n2246), .Y(n6487) );
  NAND2X1 U4277 ( .A(ram[2050]), .B(n12907), .Y(n2246) );
  OAI21X1 U4278 ( .A(n12761), .B(n12907), .C(n2247), .Y(n6488) );
  NAND2X1 U4279 ( .A(ram[2051]), .B(n12907), .Y(n2247) );
  OAI21X1 U4280 ( .A(n12755), .B(n12907), .C(n2248), .Y(n6489) );
  NAND2X1 U4281 ( .A(ram[2052]), .B(n12907), .Y(n2248) );
  OAI21X1 U4282 ( .A(n12749), .B(n12907), .C(n2249), .Y(n6490) );
  NAND2X1 U4283 ( .A(ram[2053]), .B(n12907), .Y(n2249) );
  OAI21X1 U4284 ( .A(n12743), .B(n12907), .C(n2250), .Y(n6491) );
  NAND2X1 U4285 ( .A(ram[2054]), .B(n12907), .Y(n2250) );
  OAI21X1 U4286 ( .A(n12737), .B(n12907), .C(n2251), .Y(n6492) );
  NAND2X1 U4287 ( .A(ram[2055]), .B(n12907), .Y(n2251) );
  OAI21X1 U4288 ( .A(n12731), .B(n12907), .C(n2252), .Y(n6493) );
  NAND2X1 U4289 ( .A(ram[2056]), .B(n12907), .Y(n2252) );
  OAI21X1 U4290 ( .A(n12725), .B(n12907), .C(n2253), .Y(n6494) );
  NAND2X1 U4291 ( .A(ram[2057]), .B(n12907), .Y(n2253) );
  OAI21X1 U4292 ( .A(n12719), .B(n12907), .C(n2254), .Y(n6495) );
  NAND2X1 U4293 ( .A(ram[2058]), .B(n12907), .Y(n2254) );
  OAI21X1 U4294 ( .A(n12713), .B(n12907), .C(n2255), .Y(n6496) );
  NAND2X1 U4295 ( .A(ram[2059]), .B(n12907), .Y(n2255) );
  OAI21X1 U4296 ( .A(n12707), .B(n12907), .C(n2256), .Y(n6497) );
  NAND2X1 U4297 ( .A(ram[2060]), .B(n12907), .Y(n2256) );
  OAI21X1 U4298 ( .A(n12701), .B(n12907), .C(n2257), .Y(n6498) );
  NAND2X1 U4299 ( .A(ram[2061]), .B(n12907), .Y(n2257) );
  OAI21X1 U4300 ( .A(n12693), .B(n12907), .C(n2258), .Y(n6499) );
  NAND2X1 U4301 ( .A(ram[2062]), .B(n12907), .Y(n2258) );
  OAI21X1 U4302 ( .A(n12687), .B(n12907), .C(n2259), .Y(n6500) );
  NAND2X1 U4303 ( .A(ram[2063]), .B(n12907), .Y(n2259) );
  OAI21X1 U4305 ( .A(n12777), .B(n12906), .C(n2261), .Y(n6501) );
  NAND2X1 U4306 ( .A(ram[2064]), .B(n12906), .Y(n2261) );
  OAI21X1 U4307 ( .A(n12771), .B(n12906), .C(n2262), .Y(n6502) );
  NAND2X1 U4308 ( .A(ram[2065]), .B(n12906), .Y(n2262) );
  OAI21X1 U4309 ( .A(n12766), .B(n12906), .C(n2263), .Y(n6503) );
  NAND2X1 U4310 ( .A(ram[2066]), .B(n12906), .Y(n2263) );
  OAI21X1 U4311 ( .A(n12760), .B(n12906), .C(n2264), .Y(n6504) );
  NAND2X1 U4312 ( .A(ram[2067]), .B(n12906), .Y(n2264) );
  OAI21X1 U4313 ( .A(n12754), .B(n12906), .C(n2265), .Y(n6505) );
  NAND2X1 U4314 ( .A(ram[2068]), .B(n12906), .Y(n2265) );
  OAI21X1 U4315 ( .A(n12748), .B(n12906), .C(n2266), .Y(n6506) );
  NAND2X1 U4316 ( .A(ram[2069]), .B(n12906), .Y(n2266) );
  OAI21X1 U4317 ( .A(n12742), .B(n12906), .C(n2267), .Y(n6507) );
  NAND2X1 U4318 ( .A(ram[2070]), .B(n12906), .Y(n2267) );
  OAI21X1 U4319 ( .A(n12736), .B(n12906), .C(n2268), .Y(n6508) );
  NAND2X1 U4320 ( .A(ram[2071]), .B(n12906), .Y(n2268) );
  OAI21X1 U4321 ( .A(n12730), .B(n12906), .C(n2269), .Y(n6509) );
  NAND2X1 U4322 ( .A(ram[2072]), .B(n12906), .Y(n2269) );
  OAI21X1 U4323 ( .A(n12724), .B(n12906), .C(n2270), .Y(n6510) );
  NAND2X1 U4324 ( .A(ram[2073]), .B(n12906), .Y(n2270) );
  OAI21X1 U4325 ( .A(n12718), .B(n12906), .C(n2271), .Y(n6511) );
  NAND2X1 U4326 ( .A(ram[2074]), .B(n12906), .Y(n2271) );
  OAI21X1 U4327 ( .A(n12712), .B(n12906), .C(n2272), .Y(n6512) );
  NAND2X1 U4328 ( .A(ram[2075]), .B(n12906), .Y(n2272) );
  OAI21X1 U4329 ( .A(n12706), .B(n12906), .C(n2273), .Y(n6513) );
  NAND2X1 U4330 ( .A(ram[2076]), .B(n12906), .Y(n2273) );
  OAI21X1 U4331 ( .A(n12700), .B(n12906), .C(n2274), .Y(n6514) );
  NAND2X1 U4332 ( .A(ram[2077]), .B(n12906), .Y(n2274) );
  OAI21X1 U4333 ( .A(n12693), .B(n12906), .C(n2275), .Y(n6515) );
  NAND2X1 U4334 ( .A(ram[2078]), .B(n12906), .Y(n2275) );
  OAI21X1 U4335 ( .A(n12687), .B(n12906), .C(n2276), .Y(n6516) );
  NAND2X1 U4336 ( .A(ram[2079]), .B(n12906), .Y(n2276) );
  OAI21X1 U4338 ( .A(n12775), .B(n12905), .C(n2278), .Y(n6517) );
  NAND2X1 U4339 ( .A(ram[2080]), .B(n12905), .Y(n2278) );
  OAI21X1 U4340 ( .A(n12769), .B(n12905), .C(n2279), .Y(n6518) );
  NAND2X1 U4341 ( .A(ram[2081]), .B(n12905), .Y(n2279) );
  OAI21X1 U4342 ( .A(n12762), .B(n12905), .C(n2280), .Y(n6519) );
  NAND2X1 U4343 ( .A(ram[2082]), .B(n12905), .Y(n2280) );
  OAI21X1 U4344 ( .A(n12756), .B(n12905), .C(n2281), .Y(n6520) );
  NAND2X1 U4345 ( .A(ram[2083]), .B(n12905), .Y(n2281) );
  OAI21X1 U4346 ( .A(n12750), .B(n12905), .C(n2282), .Y(n6521) );
  NAND2X1 U4347 ( .A(ram[2084]), .B(n12905), .Y(n2282) );
  OAI21X1 U4348 ( .A(n12744), .B(n12905), .C(n2283), .Y(n6522) );
  NAND2X1 U4349 ( .A(ram[2085]), .B(n12905), .Y(n2283) );
  OAI21X1 U4350 ( .A(n12738), .B(n12905), .C(n2284), .Y(n6523) );
  NAND2X1 U4351 ( .A(ram[2086]), .B(n12905), .Y(n2284) );
  OAI21X1 U4352 ( .A(n12732), .B(n12905), .C(n2285), .Y(n6524) );
  NAND2X1 U4353 ( .A(ram[2087]), .B(n12905), .Y(n2285) );
  OAI21X1 U4354 ( .A(n12726), .B(n12905), .C(n2286), .Y(n6525) );
  NAND2X1 U4355 ( .A(ram[2088]), .B(n12905), .Y(n2286) );
  OAI21X1 U4356 ( .A(n12720), .B(n12905), .C(n2287), .Y(n6526) );
  NAND2X1 U4357 ( .A(ram[2089]), .B(n12905), .Y(n2287) );
  OAI21X1 U4358 ( .A(n12714), .B(n12905), .C(n2288), .Y(n6527) );
  NAND2X1 U4359 ( .A(ram[2090]), .B(n12905), .Y(n2288) );
  OAI21X1 U4360 ( .A(n12708), .B(n12905), .C(n2289), .Y(n6528) );
  NAND2X1 U4361 ( .A(ram[2091]), .B(n12905), .Y(n2289) );
  OAI21X1 U4362 ( .A(n12702), .B(n12905), .C(n2290), .Y(n6529) );
  NAND2X1 U4363 ( .A(ram[2092]), .B(n12905), .Y(n2290) );
  OAI21X1 U4364 ( .A(n12696), .B(n12905), .C(n2291), .Y(n6530) );
  NAND2X1 U4365 ( .A(ram[2093]), .B(n12905), .Y(n2291) );
  OAI21X1 U4366 ( .A(n12691), .B(n12905), .C(n2292), .Y(n6531) );
  NAND2X1 U4367 ( .A(ram[2094]), .B(n12905), .Y(n2292) );
  OAI21X1 U4368 ( .A(n12685), .B(n12905), .C(n2293), .Y(n6532) );
  NAND2X1 U4369 ( .A(ram[2095]), .B(n12905), .Y(n2293) );
  OAI21X1 U4371 ( .A(n12774), .B(n12904), .C(n2295), .Y(n6533) );
  NAND2X1 U4372 ( .A(ram[2096]), .B(n12904), .Y(n2295) );
  OAI21X1 U4373 ( .A(n12768), .B(n12904), .C(n2296), .Y(n6534) );
  NAND2X1 U4374 ( .A(ram[2097]), .B(n12904), .Y(n2296) );
  OAI21X1 U4375 ( .A(n12763), .B(n12904), .C(n2297), .Y(n6535) );
  NAND2X1 U4376 ( .A(ram[2098]), .B(n12904), .Y(n2297) );
  OAI21X1 U4377 ( .A(n12757), .B(n12904), .C(n2298), .Y(n6536) );
  NAND2X1 U4378 ( .A(ram[2099]), .B(n12904), .Y(n2298) );
  OAI21X1 U4379 ( .A(n12751), .B(n12904), .C(n2299), .Y(n6537) );
  NAND2X1 U4380 ( .A(ram[2100]), .B(n12904), .Y(n2299) );
  OAI21X1 U4381 ( .A(n12745), .B(n12904), .C(n2300), .Y(n6538) );
  NAND2X1 U4382 ( .A(ram[2101]), .B(n12904), .Y(n2300) );
  OAI21X1 U4383 ( .A(n12739), .B(n12904), .C(n2301), .Y(n6539) );
  NAND2X1 U4384 ( .A(ram[2102]), .B(n12904), .Y(n2301) );
  OAI21X1 U4385 ( .A(n12733), .B(n12904), .C(n2302), .Y(n6540) );
  NAND2X1 U4386 ( .A(ram[2103]), .B(n12904), .Y(n2302) );
  OAI21X1 U4387 ( .A(n12727), .B(n12904), .C(n2303), .Y(n6541) );
  NAND2X1 U4388 ( .A(ram[2104]), .B(n12904), .Y(n2303) );
  OAI21X1 U4389 ( .A(n12721), .B(n12904), .C(n2304), .Y(n6542) );
  NAND2X1 U4390 ( .A(ram[2105]), .B(n12904), .Y(n2304) );
  OAI21X1 U4391 ( .A(n12715), .B(n12904), .C(n2305), .Y(n6543) );
  NAND2X1 U4392 ( .A(ram[2106]), .B(n12904), .Y(n2305) );
  OAI21X1 U4393 ( .A(n12709), .B(n12904), .C(n2306), .Y(n6544) );
  NAND2X1 U4394 ( .A(ram[2107]), .B(n12904), .Y(n2306) );
  OAI21X1 U4395 ( .A(n12703), .B(n12904), .C(n2307), .Y(n6545) );
  NAND2X1 U4396 ( .A(ram[2108]), .B(n12904), .Y(n2307) );
  OAI21X1 U4397 ( .A(n12697), .B(n12904), .C(n2308), .Y(n6546) );
  NAND2X1 U4398 ( .A(ram[2109]), .B(n12904), .Y(n2308) );
  OAI21X1 U4399 ( .A(n12690), .B(n12904), .C(n2309), .Y(n6547) );
  NAND2X1 U4400 ( .A(ram[2110]), .B(n12904), .Y(n2309) );
  OAI21X1 U4401 ( .A(n12684), .B(n12904), .C(n2310), .Y(n6548) );
  NAND2X1 U4402 ( .A(ram[2111]), .B(n12904), .Y(n2310) );
  OAI21X1 U4404 ( .A(n12778), .B(n12903), .C(n2312), .Y(n6549) );
  NAND2X1 U4405 ( .A(ram[2112]), .B(n12903), .Y(n2312) );
  OAI21X1 U4406 ( .A(n12772), .B(n12903), .C(n2313), .Y(n6550) );
  NAND2X1 U4407 ( .A(ram[2113]), .B(n12903), .Y(n2313) );
  OAI21X1 U4408 ( .A(n12763), .B(n12903), .C(n2314), .Y(n6551) );
  NAND2X1 U4409 ( .A(ram[2114]), .B(n12903), .Y(n2314) );
  OAI21X1 U4410 ( .A(n12757), .B(n12903), .C(n2315), .Y(n6552) );
  NAND2X1 U4411 ( .A(ram[2115]), .B(n12903), .Y(n2315) );
  OAI21X1 U4412 ( .A(n12751), .B(n12903), .C(n2316), .Y(n6553) );
  NAND2X1 U4413 ( .A(ram[2116]), .B(n12903), .Y(n2316) );
  OAI21X1 U4414 ( .A(n12745), .B(n12903), .C(n2317), .Y(n6554) );
  NAND2X1 U4415 ( .A(ram[2117]), .B(n12903), .Y(n2317) );
  OAI21X1 U4416 ( .A(n12739), .B(n12903), .C(n2318), .Y(n6555) );
  NAND2X1 U4417 ( .A(ram[2118]), .B(n12903), .Y(n2318) );
  OAI21X1 U4418 ( .A(n12733), .B(n12903), .C(n2319), .Y(n6556) );
  NAND2X1 U4419 ( .A(ram[2119]), .B(n12903), .Y(n2319) );
  OAI21X1 U4420 ( .A(n12727), .B(n12903), .C(n2320), .Y(n6557) );
  NAND2X1 U4421 ( .A(ram[2120]), .B(n12903), .Y(n2320) );
  OAI21X1 U4422 ( .A(n12721), .B(n12903), .C(n2321), .Y(n6558) );
  NAND2X1 U4423 ( .A(ram[2121]), .B(n12903), .Y(n2321) );
  OAI21X1 U4424 ( .A(n12715), .B(n12903), .C(n2322), .Y(n6559) );
  NAND2X1 U4425 ( .A(ram[2122]), .B(n12903), .Y(n2322) );
  OAI21X1 U4426 ( .A(n12709), .B(n12903), .C(n2323), .Y(n6560) );
  NAND2X1 U4427 ( .A(ram[2123]), .B(n12903), .Y(n2323) );
  OAI21X1 U4428 ( .A(n12703), .B(n12903), .C(n2324), .Y(n6561) );
  NAND2X1 U4429 ( .A(ram[2124]), .B(n12903), .Y(n2324) );
  OAI21X1 U4430 ( .A(n12697), .B(n12903), .C(n2325), .Y(n6562) );
  NAND2X1 U4431 ( .A(ram[2125]), .B(n12903), .Y(n2325) );
  OAI21X1 U4432 ( .A(n12694), .B(n12903), .C(n2326), .Y(n6563) );
  NAND2X1 U4433 ( .A(ram[2126]), .B(n12903), .Y(n2326) );
  OAI21X1 U4434 ( .A(n12688), .B(n12903), .C(n2327), .Y(n6564) );
  NAND2X1 U4435 ( .A(ram[2127]), .B(n12903), .Y(n2327) );
  OAI21X1 U4437 ( .A(n12779), .B(n12902), .C(n2329), .Y(n6565) );
  NAND2X1 U4438 ( .A(ram[2128]), .B(n12902), .Y(n2329) );
  OAI21X1 U4439 ( .A(n12773), .B(n12902), .C(n2330), .Y(n6566) );
  NAND2X1 U4440 ( .A(ram[2129]), .B(n12902), .Y(n2330) );
  OAI21X1 U4441 ( .A(n12762), .B(n12902), .C(n2331), .Y(n6567) );
  NAND2X1 U4442 ( .A(ram[2130]), .B(n12902), .Y(n2331) );
  OAI21X1 U4443 ( .A(n12756), .B(n12902), .C(n2332), .Y(n6568) );
  NAND2X1 U4444 ( .A(ram[2131]), .B(n12902), .Y(n2332) );
  OAI21X1 U4445 ( .A(n12750), .B(n12902), .C(n2333), .Y(n6569) );
  NAND2X1 U4446 ( .A(ram[2132]), .B(n12902), .Y(n2333) );
  OAI21X1 U4447 ( .A(n12744), .B(n12902), .C(n2334), .Y(n6570) );
  NAND2X1 U4448 ( .A(ram[2133]), .B(n12902), .Y(n2334) );
  OAI21X1 U4449 ( .A(n12738), .B(n12902), .C(n2335), .Y(n6571) );
  NAND2X1 U4450 ( .A(ram[2134]), .B(n12902), .Y(n2335) );
  OAI21X1 U4451 ( .A(n12732), .B(n12902), .C(n2336), .Y(n6572) );
  NAND2X1 U4452 ( .A(ram[2135]), .B(n12902), .Y(n2336) );
  OAI21X1 U4453 ( .A(n12726), .B(n12902), .C(n2337), .Y(n6573) );
  NAND2X1 U4454 ( .A(ram[2136]), .B(n12902), .Y(n2337) );
  OAI21X1 U4455 ( .A(n12720), .B(n12902), .C(n2338), .Y(n6574) );
  NAND2X1 U4456 ( .A(ram[2137]), .B(n12902), .Y(n2338) );
  OAI21X1 U4457 ( .A(n12714), .B(n12902), .C(n2339), .Y(n6575) );
  NAND2X1 U4458 ( .A(ram[2138]), .B(n12902), .Y(n2339) );
  OAI21X1 U4459 ( .A(n12708), .B(n12902), .C(n2340), .Y(n6576) );
  NAND2X1 U4460 ( .A(ram[2139]), .B(n12902), .Y(n2340) );
  OAI21X1 U4461 ( .A(n12702), .B(n12902), .C(n2341), .Y(n6577) );
  NAND2X1 U4462 ( .A(ram[2140]), .B(n12902), .Y(n2341) );
  OAI21X1 U4463 ( .A(n12696), .B(n12902), .C(n2342), .Y(n6578) );
  NAND2X1 U4464 ( .A(ram[2141]), .B(n12902), .Y(n2342) );
  OAI21X1 U4465 ( .A(n12695), .B(n12902), .C(n2343), .Y(n6579) );
  NAND2X1 U4466 ( .A(ram[2142]), .B(n12902), .Y(n2343) );
  OAI21X1 U4467 ( .A(n12689), .B(n12902), .C(n2344), .Y(n6580) );
  NAND2X1 U4468 ( .A(ram[2143]), .B(n12902), .Y(n2344) );
  OAI21X1 U4470 ( .A(n12779), .B(n12901), .C(n2346), .Y(n6581) );
  NAND2X1 U4471 ( .A(ram[2144]), .B(n12901), .Y(n2346) );
  OAI21X1 U4472 ( .A(n12773), .B(n12901), .C(n2347), .Y(n6582) );
  NAND2X1 U4473 ( .A(ram[2145]), .B(n12901), .Y(n2347) );
  OAI21X1 U4474 ( .A(n12767), .B(n12901), .C(n2348), .Y(n6583) );
  NAND2X1 U4475 ( .A(ram[2146]), .B(n12901), .Y(n2348) );
  OAI21X1 U4476 ( .A(n12761), .B(n12901), .C(n2349), .Y(n6584) );
  NAND2X1 U4477 ( .A(ram[2147]), .B(n12901), .Y(n2349) );
  OAI21X1 U4478 ( .A(n12755), .B(n12901), .C(n2350), .Y(n6585) );
  NAND2X1 U4479 ( .A(ram[2148]), .B(n12901), .Y(n2350) );
  OAI21X1 U4480 ( .A(n12749), .B(n12901), .C(n2351), .Y(n6586) );
  NAND2X1 U4481 ( .A(ram[2149]), .B(n12901), .Y(n2351) );
  OAI21X1 U4482 ( .A(n12743), .B(n12901), .C(n2352), .Y(n6587) );
  NAND2X1 U4483 ( .A(ram[2150]), .B(n12901), .Y(n2352) );
  OAI21X1 U4484 ( .A(n12737), .B(n12901), .C(n2353), .Y(n6588) );
  NAND2X1 U4485 ( .A(ram[2151]), .B(n12901), .Y(n2353) );
  OAI21X1 U4486 ( .A(n12731), .B(n12901), .C(n2354), .Y(n6589) );
  NAND2X1 U4487 ( .A(ram[2152]), .B(n12901), .Y(n2354) );
  OAI21X1 U4488 ( .A(n12725), .B(n12901), .C(n2355), .Y(n6590) );
  NAND2X1 U4489 ( .A(ram[2153]), .B(n12901), .Y(n2355) );
  OAI21X1 U4490 ( .A(n12719), .B(n12901), .C(n2356), .Y(n6591) );
  NAND2X1 U4491 ( .A(ram[2154]), .B(n12901), .Y(n2356) );
  OAI21X1 U4492 ( .A(n12713), .B(n12901), .C(n2357), .Y(n6592) );
  NAND2X1 U4493 ( .A(ram[2155]), .B(n12901), .Y(n2357) );
  OAI21X1 U4494 ( .A(n12707), .B(n12901), .C(n2358), .Y(n6593) );
  NAND2X1 U4495 ( .A(ram[2156]), .B(n12901), .Y(n2358) );
  OAI21X1 U4496 ( .A(n12701), .B(n12901), .C(n2359), .Y(n6594) );
  NAND2X1 U4497 ( .A(ram[2157]), .B(n12901), .Y(n2359) );
  OAI21X1 U4498 ( .A(n12695), .B(n12901), .C(n2360), .Y(n6595) );
  NAND2X1 U4499 ( .A(ram[2158]), .B(n12901), .Y(n2360) );
  OAI21X1 U4500 ( .A(n12689), .B(n12901), .C(n2361), .Y(n6596) );
  NAND2X1 U4501 ( .A(ram[2159]), .B(n12901), .Y(n2361) );
  OAI21X1 U4503 ( .A(n12778), .B(n12900), .C(n2363), .Y(n6597) );
  NAND2X1 U4504 ( .A(ram[2160]), .B(n12900), .Y(n2363) );
  OAI21X1 U4505 ( .A(n12772), .B(n12900), .C(n2364), .Y(n6598) );
  NAND2X1 U4506 ( .A(ram[2161]), .B(n12900), .Y(n2364) );
  OAI21X1 U4507 ( .A(n12766), .B(n12900), .C(n2365), .Y(n6599) );
  NAND2X1 U4508 ( .A(ram[2162]), .B(n12900), .Y(n2365) );
  OAI21X1 U4509 ( .A(n12760), .B(n12900), .C(n2366), .Y(n6600) );
  NAND2X1 U4510 ( .A(ram[2163]), .B(n12900), .Y(n2366) );
  OAI21X1 U4511 ( .A(n12754), .B(n12900), .C(n2367), .Y(n6601) );
  NAND2X1 U4512 ( .A(ram[2164]), .B(n12900), .Y(n2367) );
  OAI21X1 U4513 ( .A(n12748), .B(n12900), .C(n2368), .Y(n6602) );
  NAND2X1 U4514 ( .A(ram[2165]), .B(n12900), .Y(n2368) );
  OAI21X1 U4515 ( .A(n12742), .B(n12900), .C(n2369), .Y(n6603) );
  NAND2X1 U4516 ( .A(ram[2166]), .B(n12900), .Y(n2369) );
  OAI21X1 U4517 ( .A(n12736), .B(n12900), .C(n2370), .Y(n6604) );
  NAND2X1 U4518 ( .A(ram[2167]), .B(n12900), .Y(n2370) );
  OAI21X1 U4519 ( .A(n12730), .B(n12900), .C(n2371), .Y(n6605) );
  NAND2X1 U4520 ( .A(ram[2168]), .B(n12900), .Y(n2371) );
  OAI21X1 U4521 ( .A(n12724), .B(n12900), .C(n2372), .Y(n6606) );
  NAND2X1 U4522 ( .A(ram[2169]), .B(n12900), .Y(n2372) );
  OAI21X1 U4523 ( .A(n12718), .B(n12900), .C(n2373), .Y(n6607) );
  NAND2X1 U4524 ( .A(ram[2170]), .B(n12900), .Y(n2373) );
  OAI21X1 U4525 ( .A(n12712), .B(n12900), .C(n2374), .Y(n6608) );
  NAND2X1 U4526 ( .A(ram[2171]), .B(n12900), .Y(n2374) );
  OAI21X1 U4527 ( .A(n12706), .B(n12900), .C(n2375), .Y(n6609) );
  NAND2X1 U4528 ( .A(ram[2172]), .B(n12900), .Y(n2375) );
  OAI21X1 U4529 ( .A(n12700), .B(n12900), .C(n2376), .Y(n6610) );
  NAND2X1 U4530 ( .A(ram[2173]), .B(n12900), .Y(n2376) );
  OAI21X1 U4531 ( .A(n12694), .B(n12900), .C(n2377), .Y(n6611) );
  NAND2X1 U4532 ( .A(ram[2174]), .B(n12900), .Y(n2377) );
  OAI21X1 U4533 ( .A(n12688), .B(n12900), .C(n2378), .Y(n6612) );
  NAND2X1 U4534 ( .A(ram[2175]), .B(n12900), .Y(n2378) );
  OAI21X1 U4536 ( .A(n12777), .B(n12899), .C(n2380), .Y(n6613) );
  NAND2X1 U4537 ( .A(ram[2176]), .B(n12899), .Y(n2380) );
  OAI21X1 U4538 ( .A(n12771), .B(n12899), .C(n2381), .Y(n6614) );
  NAND2X1 U4539 ( .A(ram[2177]), .B(n12899), .Y(n2381) );
  OAI21X1 U4540 ( .A(n12765), .B(n12899), .C(n2382), .Y(n6615) );
  NAND2X1 U4541 ( .A(ram[2178]), .B(n12899), .Y(n2382) );
  OAI21X1 U4542 ( .A(n12759), .B(n12899), .C(n2383), .Y(n6616) );
  NAND2X1 U4543 ( .A(ram[2179]), .B(n12899), .Y(n2383) );
  OAI21X1 U4544 ( .A(n12753), .B(n12899), .C(n2384), .Y(n6617) );
  NAND2X1 U4545 ( .A(ram[2180]), .B(n12899), .Y(n2384) );
  OAI21X1 U4546 ( .A(n12747), .B(n12899), .C(n2385), .Y(n6618) );
  NAND2X1 U4547 ( .A(ram[2181]), .B(n12899), .Y(n2385) );
  OAI21X1 U4548 ( .A(n12741), .B(n12899), .C(n2386), .Y(n6619) );
  NAND2X1 U4549 ( .A(ram[2182]), .B(n12899), .Y(n2386) );
  OAI21X1 U4550 ( .A(n12735), .B(n12899), .C(n2387), .Y(n6620) );
  NAND2X1 U4551 ( .A(ram[2183]), .B(n12899), .Y(n2387) );
  OAI21X1 U4552 ( .A(n12729), .B(n12899), .C(n2388), .Y(n6621) );
  NAND2X1 U4553 ( .A(ram[2184]), .B(n12899), .Y(n2388) );
  OAI21X1 U4554 ( .A(n12723), .B(n12899), .C(n2389), .Y(n6622) );
  NAND2X1 U4555 ( .A(ram[2185]), .B(n12899), .Y(n2389) );
  OAI21X1 U4556 ( .A(n12717), .B(n12899), .C(n2390), .Y(n6623) );
  NAND2X1 U4557 ( .A(ram[2186]), .B(n12899), .Y(n2390) );
  OAI21X1 U4558 ( .A(n12711), .B(n12899), .C(n2391), .Y(n6624) );
  NAND2X1 U4559 ( .A(ram[2187]), .B(n12899), .Y(n2391) );
  OAI21X1 U4560 ( .A(n12705), .B(n12899), .C(n2392), .Y(n6625) );
  NAND2X1 U4561 ( .A(ram[2188]), .B(n12899), .Y(n2392) );
  OAI21X1 U4562 ( .A(n12699), .B(n12899), .C(n2393), .Y(n6626) );
  NAND2X1 U4563 ( .A(ram[2189]), .B(n12899), .Y(n2393) );
  OAI21X1 U4564 ( .A(n12693), .B(n12899), .C(n2394), .Y(n6627) );
  NAND2X1 U4565 ( .A(ram[2190]), .B(n12899), .Y(n2394) );
  OAI21X1 U4566 ( .A(n12687), .B(n12899), .C(n2395), .Y(n6628) );
  NAND2X1 U4567 ( .A(ram[2191]), .B(n12899), .Y(n2395) );
  OAI21X1 U4569 ( .A(n12778), .B(n12898), .C(n2397), .Y(n6629) );
  NAND2X1 U4570 ( .A(ram[2192]), .B(n12898), .Y(n2397) );
  OAI21X1 U4571 ( .A(n12772), .B(n12898), .C(n2398), .Y(n6630) );
  NAND2X1 U4572 ( .A(ram[2193]), .B(n12898), .Y(n2398) );
  OAI21X1 U4573 ( .A(n12763), .B(n12898), .C(n2399), .Y(n6631) );
  NAND2X1 U4574 ( .A(ram[2194]), .B(n12898), .Y(n2399) );
  OAI21X1 U4575 ( .A(n12757), .B(n12898), .C(n2400), .Y(n6632) );
  NAND2X1 U4576 ( .A(ram[2195]), .B(n12898), .Y(n2400) );
  OAI21X1 U4577 ( .A(n12751), .B(n12898), .C(n2401), .Y(n6633) );
  NAND2X1 U4578 ( .A(ram[2196]), .B(n12898), .Y(n2401) );
  OAI21X1 U4579 ( .A(n12745), .B(n12898), .C(n2402), .Y(n6634) );
  NAND2X1 U4580 ( .A(ram[2197]), .B(n12898), .Y(n2402) );
  OAI21X1 U4581 ( .A(n12739), .B(n12898), .C(n2403), .Y(n6635) );
  NAND2X1 U4582 ( .A(ram[2198]), .B(n12898), .Y(n2403) );
  OAI21X1 U4583 ( .A(n12733), .B(n12898), .C(n2404), .Y(n6636) );
  NAND2X1 U4584 ( .A(ram[2199]), .B(n12898), .Y(n2404) );
  OAI21X1 U4585 ( .A(n12727), .B(n12898), .C(n2405), .Y(n6637) );
  NAND2X1 U4586 ( .A(ram[2200]), .B(n12898), .Y(n2405) );
  OAI21X1 U4587 ( .A(n12721), .B(n12898), .C(n2406), .Y(n6638) );
  NAND2X1 U4588 ( .A(ram[2201]), .B(n12898), .Y(n2406) );
  OAI21X1 U4589 ( .A(n12715), .B(n12898), .C(n2407), .Y(n6639) );
  NAND2X1 U4590 ( .A(ram[2202]), .B(n12898), .Y(n2407) );
  OAI21X1 U4591 ( .A(n12709), .B(n12898), .C(n2408), .Y(n6640) );
  NAND2X1 U4592 ( .A(ram[2203]), .B(n12898), .Y(n2408) );
  OAI21X1 U4593 ( .A(n12703), .B(n12898), .C(n2409), .Y(n6641) );
  NAND2X1 U4594 ( .A(ram[2204]), .B(n12898), .Y(n2409) );
  OAI21X1 U4595 ( .A(n12697), .B(n12898), .C(n2410), .Y(n6642) );
  NAND2X1 U4596 ( .A(ram[2205]), .B(n12898), .Y(n2410) );
  OAI21X1 U4597 ( .A(n12694), .B(n12898), .C(n2411), .Y(n6643) );
  NAND2X1 U4598 ( .A(ram[2206]), .B(n12898), .Y(n2411) );
  OAI21X1 U4599 ( .A(n12688), .B(n12898), .C(n2412), .Y(n6644) );
  NAND2X1 U4600 ( .A(ram[2207]), .B(n12898), .Y(n2412) );
  OAI21X1 U4602 ( .A(n12775), .B(n12897), .C(n2414), .Y(n6645) );
  NAND2X1 U4603 ( .A(ram[2208]), .B(n12897), .Y(n2414) );
  OAI21X1 U4604 ( .A(n12769), .B(n12897), .C(n2415), .Y(n6646) );
  NAND2X1 U4605 ( .A(ram[2209]), .B(n12897), .Y(n2415) );
  OAI21X1 U4606 ( .A(n12765), .B(n12897), .C(n2416), .Y(n6647) );
  NAND2X1 U4607 ( .A(ram[2210]), .B(n12897), .Y(n2416) );
  OAI21X1 U4608 ( .A(n12759), .B(n12897), .C(n2417), .Y(n6648) );
  NAND2X1 U4609 ( .A(ram[2211]), .B(n12897), .Y(n2417) );
  OAI21X1 U4610 ( .A(n12753), .B(n12897), .C(n2418), .Y(n6649) );
  NAND2X1 U4611 ( .A(ram[2212]), .B(n12897), .Y(n2418) );
  OAI21X1 U4612 ( .A(n12747), .B(n12897), .C(n2419), .Y(n6650) );
  NAND2X1 U4613 ( .A(ram[2213]), .B(n12897), .Y(n2419) );
  OAI21X1 U4614 ( .A(n12741), .B(n12897), .C(n2420), .Y(n6651) );
  NAND2X1 U4615 ( .A(ram[2214]), .B(n12897), .Y(n2420) );
  OAI21X1 U4616 ( .A(n12735), .B(n12897), .C(n2421), .Y(n6652) );
  NAND2X1 U4617 ( .A(ram[2215]), .B(n12897), .Y(n2421) );
  OAI21X1 U4618 ( .A(n12729), .B(n12897), .C(n2422), .Y(n6653) );
  NAND2X1 U4619 ( .A(ram[2216]), .B(n12897), .Y(n2422) );
  OAI21X1 U4620 ( .A(n12723), .B(n12897), .C(n2423), .Y(n6654) );
  NAND2X1 U4621 ( .A(ram[2217]), .B(n12897), .Y(n2423) );
  OAI21X1 U4622 ( .A(n12717), .B(n12897), .C(n2424), .Y(n6655) );
  NAND2X1 U4623 ( .A(ram[2218]), .B(n12897), .Y(n2424) );
  OAI21X1 U4624 ( .A(n12711), .B(n12897), .C(n2425), .Y(n6656) );
  NAND2X1 U4625 ( .A(ram[2219]), .B(n12897), .Y(n2425) );
  OAI21X1 U4626 ( .A(n12705), .B(n12897), .C(n2426), .Y(n6657) );
  NAND2X1 U4627 ( .A(ram[2220]), .B(n12897), .Y(n2426) );
  OAI21X1 U4628 ( .A(n12699), .B(n12897), .C(n2427), .Y(n6658) );
  NAND2X1 U4629 ( .A(ram[2221]), .B(n12897), .Y(n2427) );
  OAI21X1 U4630 ( .A(n12691), .B(n12897), .C(n2428), .Y(n6659) );
  NAND2X1 U4631 ( .A(ram[2222]), .B(n12897), .Y(n2428) );
  OAI21X1 U4632 ( .A(n12685), .B(n12897), .C(n2429), .Y(n6660) );
  NAND2X1 U4633 ( .A(ram[2223]), .B(n12897), .Y(n2429) );
  OAI21X1 U4635 ( .A(n12774), .B(n12896), .C(n2431), .Y(n6661) );
  NAND2X1 U4636 ( .A(ram[2224]), .B(n12896), .Y(n2431) );
  OAI21X1 U4637 ( .A(n12768), .B(n12896), .C(n2432), .Y(n6662) );
  NAND2X1 U4638 ( .A(ram[2225]), .B(n12896), .Y(n2432) );
  OAI21X1 U4639 ( .A(n12765), .B(n12896), .C(n2433), .Y(n6663) );
  NAND2X1 U4640 ( .A(ram[2226]), .B(n12896), .Y(n2433) );
  OAI21X1 U4641 ( .A(n12759), .B(n12896), .C(n2434), .Y(n6664) );
  NAND2X1 U4642 ( .A(ram[2227]), .B(n12896), .Y(n2434) );
  OAI21X1 U4643 ( .A(n12753), .B(n12896), .C(n2435), .Y(n6665) );
  NAND2X1 U4644 ( .A(ram[2228]), .B(n12896), .Y(n2435) );
  OAI21X1 U4645 ( .A(n12747), .B(n12896), .C(n2436), .Y(n6666) );
  NAND2X1 U4646 ( .A(ram[2229]), .B(n12896), .Y(n2436) );
  OAI21X1 U4647 ( .A(n12741), .B(n12896), .C(n2437), .Y(n6667) );
  NAND2X1 U4648 ( .A(ram[2230]), .B(n12896), .Y(n2437) );
  OAI21X1 U4649 ( .A(n12735), .B(n12896), .C(n2438), .Y(n6668) );
  NAND2X1 U4650 ( .A(ram[2231]), .B(n12896), .Y(n2438) );
  OAI21X1 U4651 ( .A(n12729), .B(n12896), .C(n2439), .Y(n6669) );
  NAND2X1 U4652 ( .A(ram[2232]), .B(n12896), .Y(n2439) );
  OAI21X1 U4653 ( .A(n12723), .B(n12896), .C(n2440), .Y(n6670) );
  NAND2X1 U4654 ( .A(ram[2233]), .B(n12896), .Y(n2440) );
  OAI21X1 U4655 ( .A(n12717), .B(n12896), .C(n2441), .Y(n6671) );
  NAND2X1 U4656 ( .A(ram[2234]), .B(n12896), .Y(n2441) );
  OAI21X1 U4657 ( .A(n12711), .B(n12896), .C(n2442), .Y(n6672) );
  NAND2X1 U4658 ( .A(ram[2235]), .B(n12896), .Y(n2442) );
  OAI21X1 U4659 ( .A(n12705), .B(n12896), .C(n2443), .Y(n6673) );
  NAND2X1 U4660 ( .A(ram[2236]), .B(n12896), .Y(n2443) );
  OAI21X1 U4661 ( .A(n12699), .B(n12896), .C(n2444), .Y(n6674) );
  NAND2X1 U4662 ( .A(ram[2237]), .B(n12896), .Y(n2444) );
  OAI21X1 U4663 ( .A(n12690), .B(n12896), .C(n2445), .Y(n6675) );
  NAND2X1 U4664 ( .A(ram[2238]), .B(n12896), .Y(n2445) );
  OAI21X1 U4665 ( .A(n12684), .B(n12896), .C(n2446), .Y(n6676) );
  NAND2X1 U4666 ( .A(ram[2239]), .B(n12896), .Y(n2446) );
  OAI21X1 U4668 ( .A(n12776), .B(n12895), .C(n2448), .Y(n6677) );
  NAND2X1 U4669 ( .A(ram[2240]), .B(n12895), .Y(n2448) );
  OAI21X1 U4670 ( .A(n12770), .B(n12895), .C(n2449), .Y(n6678) );
  NAND2X1 U4671 ( .A(ram[2241]), .B(n12895), .Y(n2449) );
  OAI21X1 U4672 ( .A(n12767), .B(n12895), .C(n2450), .Y(n6679) );
  NAND2X1 U4673 ( .A(ram[2242]), .B(n12895), .Y(n2450) );
  OAI21X1 U4674 ( .A(n12761), .B(n12895), .C(n2451), .Y(n6680) );
  NAND2X1 U4675 ( .A(ram[2243]), .B(n12895), .Y(n2451) );
  OAI21X1 U4676 ( .A(n12755), .B(n12895), .C(n2452), .Y(n6681) );
  NAND2X1 U4677 ( .A(ram[2244]), .B(n12895), .Y(n2452) );
  OAI21X1 U4678 ( .A(n12749), .B(n12895), .C(n2453), .Y(n6682) );
  NAND2X1 U4679 ( .A(ram[2245]), .B(n12895), .Y(n2453) );
  OAI21X1 U4680 ( .A(n12743), .B(n12895), .C(n2454), .Y(n6683) );
  NAND2X1 U4681 ( .A(ram[2246]), .B(n12895), .Y(n2454) );
  OAI21X1 U4682 ( .A(n12737), .B(n12895), .C(n2455), .Y(n6684) );
  NAND2X1 U4683 ( .A(ram[2247]), .B(n12895), .Y(n2455) );
  OAI21X1 U4684 ( .A(n12731), .B(n12895), .C(n2456), .Y(n6685) );
  NAND2X1 U4685 ( .A(ram[2248]), .B(n12895), .Y(n2456) );
  OAI21X1 U4686 ( .A(n12725), .B(n12895), .C(n2457), .Y(n6686) );
  NAND2X1 U4687 ( .A(ram[2249]), .B(n12895), .Y(n2457) );
  OAI21X1 U4688 ( .A(n12719), .B(n12895), .C(n2458), .Y(n6687) );
  NAND2X1 U4689 ( .A(ram[2250]), .B(n12895), .Y(n2458) );
  OAI21X1 U4690 ( .A(n12713), .B(n12895), .C(n2459), .Y(n6688) );
  NAND2X1 U4691 ( .A(ram[2251]), .B(n12895), .Y(n2459) );
  OAI21X1 U4692 ( .A(n12707), .B(n12895), .C(n2460), .Y(n6689) );
  NAND2X1 U4693 ( .A(ram[2252]), .B(n12895), .Y(n2460) );
  OAI21X1 U4694 ( .A(n12701), .B(n12895), .C(n2461), .Y(n6690) );
  NAND2X1 U4695 ( .A(ram[2253]), .B(n12895), .Y(n2461) );
  OAI21X1 U4696 ( .A(n12692), .B(n12895), .C(n2462), .Y(n6691) );
  NAND2X1 U4697 ( .A(ram[2254]), .B(n12895), .Y(n2462) );
  OAI21X1 U4698 ( .A(n12686), .B(n12895), .C(n2463), .Y(n6692) );
  NAND2X1 U4699 ( .A(ram[2255]), .B(n12895), .Y(n2463) );
  OAI21X1 U4701 ( .A(n12775), .B(n12894), .C(n2465), .Y(n6693) );
  NAND2X1 U4702 ( .A(ram[2256]), .B(n12894), .Y(n2465) );
  OAI21X1 U4703 ( .A(n12769), .B(n12894), .C(n2466), .Y(n6694) );
  NAND2X1 U4704 ( .A(ram[2257]), .B(n12894), .Y(n2466) );
  OAI21X1 U4705 ( .A(n12764), .B(n12894), .C(n2467), .Y(n6695) );
  NAND2X1 U4706 ( .A(ram[2258]), .B(n12894), .Y(n2467) );
  OAI21X1 U4707 ( .A(n12758), .B(n12894), .C(n2468), .Y(n6696) );
  NAND2X1 U4708 ( .A(ram[2259]), .B(n12894), .Y(n2468) );
  OAI21X1 U4709 ( .A(n12752), .B(n12894), .C(n2469), .Y(n6697) );
  NAND2X1 U4710 ( .A(ram[2260]), .B(n12894), .Y(n2469) );
  OAI21X1 U4711 ( .A(n12746), .B(n12894), .C(n2470), .Y(n6698) );
  NAND2X1 U4712 ( .A(ram[2261]), .B(n12894), .Y(n2470) );
  OAI21X1 U4713 ( .A(n12740), .B(n12894), .C(n2471), .Y(n6699) );
  NAND2X1 U4714 ( .A(ram[2262]), .B(n12894), .Y(n2471) );
  OAI21X1 U4715 ( .A(n12734), .B(n12894), .C(n2472), .Y(n6700) );
  NAND2X1 U4716 ( .A(ram[2263]), .B(n12894), .Y(n2472) );
  OAI21X1 U4717 ( .A(n12728), .B(n12894), .C(n2473), .Y(n6701) );
  NAND2X1 U4718 ( .A(ram[2264]), .B(n12894), .Y(n2473) );
  OAI21X1 U4719 ( .A(n12722), .B(n12894), .C(n2474), .Y(n6702) );
  NAND2X1 U4720 ( .A(ram[2265]), .B(n12894), .Y(n2474) );
  OAI21X1 U4721 ( .A(n12716), .B(n12894), .C(n2475), .Y(n6703) );
  NAND2X1 U4722 ( .A(ram[2266]), .B(n12894), .Y(n2475) );
  OAI21X1 U4723 ( .A(n12710), .B(n12894), .C(n2476), .Y(n6704) );
  NAND2X1 U4724 ( .A(ram[2267]), .B(n12894), .Y(n2476) );
  OAI21X1 U4725 ( .A(n12704), .B(n12894), .C(n2477), .Y(n6705) );
  NAND2X1 U4726 ( .A(ram[2268]), .B(n12894), .Y(n2477) );
  OAI21X1 U4727 ( .A(n12698), .B(n12894), .C(n2478), .Y(n6706) );
  NAND2X1 U4728 ( .A(ram[2269]), .B(n12894), .Y(n2478) );
  OAI21X1 U4729 ( .A(n12691), .B(n12894), .C(n2479), .Y(n6707) );
  NAND2X1 U4730 ( .A(ram[2270]), .B(n12894), .Y(n2479) );
  OAI21X1 U4731 ( .A(n12685), .B(n12894), .C(n2480), .Y(n6708) );
  NAND2X1 U4732 ( .A(ram[2271]), .B(n12894), .Y(n2480) );
  OAI21X1 U4734 ( .A(n12775), .B(n12893), .C(n2482), .Y(n6709) );
  NAND2X1 U4735 ( .A(ram[2272]), .B(n12893), .Y(n2482) );
  OAI21X1 U4736 ( .A(n12769), .B(n12893), .C(n2483), .Y(n6710) );
  NAND2X1 U4737 ( .A(ram[2273]), .B(n12893), .Y(n2483) );
  OAI21X1 U4738 ( .A(n12762), .B(n12893), .C(n2484), .Y(n6711) );
  NAND2X1 U4739 ( .A(ram[2274]), .B(n12893), .Y(n2484) );
  OAI21X1 U4740 ( .A(n12756), .B(n12893), .C(n2485), .Y(n6712) );
  NAND2X1 U4741 ( .A(ram[2275]), .B(n12893), .Y(n2485) );
  OAI21X1 U4742 ( .A(n12750), .B(n12893), .C(n2486), .Y(n6713) );
  NAND2X1 U4743 ( .A(ram[2276]), .B(n12893), .Y(n2486) );
  OAI21X1 U4744 ( .A(n12744), .B(n12893), .C(n2487), .Y(n6714) );
  NAND2X1 U4745 ( .A(ram[2277]), .B(n12893), .Y(n2487) );
  OAI21X1 U4746 ( .A(n12738), .B(n12893), .C(n2488), .Y(n6715) );
  NAND2X1 U4747 ( .A(ram[2278]), .B(n12893), .Y(n2488) );
  OAI21X1 U4748 ( .A(n12732), .B(n12893), .C(n2489), .Y(n6716) );
  NAND2X1 U4749 ( .A(ram[2279]), .B(n12893), .Y(n2489) );
  OAI21X1 U4750 ( .A(n12726), .B(n12893), .C(n2490), .Y(n6717) );
  NAND2X1 U4751 ( .A(ram[2280]), .B(n12893), .Y(n2490) );
  OAI21X1 U4752 ( .A(n12720), .B(n12893), .C(n2491), .Y(n6718) );
  NAND2X1 U4753 ( .A(ram[2281]), .B(n12893), .Y(n2491) );
  OAI21X1 U4754 ( .A(n12714), .B(n12893), .C(n2492), .Y(n6719) );
  NAND2X1 U4755 ( .A(ram[2282]), .B(n12893), .Y(n2492) );
  OAI21X1 U4756 ( .A(n12708), .B(n12893), .C(n2493), .Y(n6720) );
  NAND2X1 U4757 ( .A(ram[2283]), .B(n12893), .Y(n2493) );
  OAI21X1 U4758 ( .A(n12702), .B(n12893), .C(n2494), .Y(n6721) );
  NAND2X1 U4759 ( .A(ram[2284]), .B(n12893), .Y(n2494) );
  OAI21X1 U4760 ( .A(n12696), .B(n12893), .C(n2495), .Y(n6722) );
  NAND2X1 U4761 ( .A(ram[2285]), .B(n12893), .Y(n2495) );
  OAI21X1 U4762 ( .A(n12691), .B(n12893), .C(n2496), .Y(n6723) );
  NAND2X1 U4763 ( .A(ram[2286]), .B(n12893), .Y(n2496) );
  OAI21X1 U4764 ( .A(n12685), .B(n12893), .C(n2497), .Y(n6724) );
  NAND2X1 U4765 ( .A(ram[2287]), .B(n12893), .Y(n2497) );
  OAI21X1 U4767 ( .A(n12779), .B(n12892), .C(n2499), .Y(n6725) );
  NAND2X1 U4768 ( .A(ram[2288]), .B(n12892), .Y(n2499) );
  OAI21X1 U4769 ( .A(n12773), .B(n12892), .C(n2500), .Y(n6726) );
  NAND2X1 U4770 ( .A(ram[2289]), .B(n12892), .Y(n2500) );
  OAI21X1 U4771 ( .A(n12762), .B(n12892), .C(n2501), .Y(n6727) );
  NAND2X1 U4772 ( .A(ram[2290]), .B(n12892), .Y(n2501) );
  OAI21X1 U4773 ( .A(n12756), .B(n12892), .C(n2502), .Y(n6728) );
  NAND2X1 U4774 ( .A(ram[2291]), .B(n12892), .Y(n2502) );
  OAI21X1 U4775 ( .A(n12750), .B(n12892), .C(n2503), .Y(n6729) );
  NAND2X1 U4776 ( .A(ram[2292]), .B(n12892), .Y(n2503) );
  OAI21X1 U4777 ( .A(n12744), .B(n12892), .C(n2504), .Y(n6730) );
  NAND2X1 U4778 ( .A(ram[2293]), .B(n12892), .Y(n2504) );
  OAI21X1 U4779 ( .A(n12738), .B(n12892), .C(n2505), .Y(n6731) );
  NAND2X1 U4780 ( .A(ram[2294]), .B(n12892), .Y(n2505) );
  OAI21X1 U4781 ( .A(n12732), .B(n12892), .C(n2506), .Y(n6732) );
  NAND2X1 U4782 ( .A(ram[2295]), .B(n12892), .Y(n2506) );
  OAI21X1 U4783 ( .A(n12726), .B(n12892), .C(n2507), .Y(n6733) );
  NAND2X1 U4784 ( .A(ram[2296]), .B(n12892), .Y(n2507) );
  OAI21X1 U4785 ( .A(n12720), .B(n12892), .C(n2508), .Y(n6734) );
  NAND2X1 U4786 ( .A(ram[2297]), .B(n12892), .Y(n2508) );
  OAI21X1 U4787 ( .A(n12714), .B(n12892), .C(n2509), .Y(n6735) );
  NAND2X1 U4788 ( .A(ram[2298]), .B(n12892), .Y(n2509) );
  OAI21X1 U4789 ( .A(n12708), .B(n12892), .C(n2510), .Y(n6736) );
  NAND2X1 U4790 ( .A(ram[2299]), .B(n12892), .Y(n2510) );
  OAI21X1 U4791 ( .A(n12702), .B(n12892), .C(n2511), .Y(n6737) );
  NAND2X1 U4792 ( .A(ram[2300]), .B(n12892), .Y(n2511) );
  OAI21X1 U4793 ( .A(n12696), .B(n12892), .C(n2512), .Y(n6738) );
  NAND2X1 U4794 ( .A(ram[2301]), .B(n12892), .Y(n2512) );
  OAI21X1 U4795 ( .A(n12695), .B(n12892), .C(n2513), .Y(n6739) );
  NAND2X1 U4796 ( .A(ram[2302]), .B(n12892), .Y(n2513) );
  OAI21X1 U4797 ( .A(n12689), .B(n12892), .C(n2514), .Y(n6740) );
  NAND2X1 U4798 ( .A(ram[2303]), .B(n12892), .Y(n2514) );
  NAND3X1 U4800 ( .A(mem_write_en), .B(n327), .C(n2516), .Y(n2515) );
  OAI21X1 U4801 ( .A(n12774), .B(n12891), .C(n2518), .Y(n6741) );
  NAND2X1 U4802 ( .A(ram[2304]), .B(n12891), .Y(n2518) );
  OAI21X1 U4803 ( .A(n12768), .B(n12891), .C(n2519), .Y(n6742) );
  NAND2X1 U4804 ( .A(ram[2305]), .B(n12891), .Y(n2519) );
  OAI21X1 U4805 ( .A(n12763), .B(n12891), .C(n2520), .Y(n6743) );
  NAND2X1 U4806 ( .A(ram[2306]), .B(n12891), .Y(n2520) );
  OAI21X1 U4807 ( .A(n12757), .B(n12891), .C(n2521), .Y(n6744) );
  NAND2X1 U4808 ( .A(ram[2307]), .B(n12891), .Y(n2521) );
  OAI21X1 U4809 ( .A(n12751), .B(n12891), .C(n2522), .Y(n6745) );
  NAND2X1 U4810 ( .A(ram[2308]), .B(n12891), .Y(n2522) );
  OAI21X1 U4811 ( .A(n12745), .B(n12891), .C(n2523), .Y(n6746) );
  NAND2X1 U4812 ( .A(ram[2309]), .B(n12891), .Y(n2523) );
  OAI21X1 U4813 ( .A(n12739), .B(n12891), .C(n2524), .Y(n6747) );
  NAND2X1 U4814 ( .A(ram[2310]), .B(n12891), .Y(n2524) );
  OAI21X1 U4815 ( .A(n12733), .B(n12891), .C(n2525), .Y(n6748) );
  NAND2X1 U4816 ( .A(ram[2311]), .B(n12891), .Y(n2525) );
  OAI21X1 U4817 ( .A(n12727), .B(n12891), .C(n2526), .Y(n6749) );
  NAND2X1 U4818 ( .A(ram[2312]), .B(n12891), .Y(n2526) );
  OAI21X1 U4819 ( .A(n12721), .B(n12891), .C(n2527), .Y(n6750) );
  NAND2X1 U4820 ( .A(ram[2313]), .B(n12891), .Y(n2527) );
  OAI21X1 U4821 ( .A(n12715), .B(n12891), .C(n2528), .Y(n6751) );
  NAND2X1 U4822 ( .A(ram[2314]), .B(n12891), .Y(n2528) );
  OAI21X1 U4823 ( .A(n12709), .B(n12891), .C(n2529), .Y(n6752) );
  NAND2X1 U4824 ( .A(ram[2315]), .B(n12891), .Y(n2529) );
  OAI21X1 U4825 ( .A(n12703), .B(n12891), .C(n2530), .Y(n6753) );
  NAND2X1 U4826 ( .A(ram[2316]), .B(n12891), .Y(n2530) );
  OAI21X1 U4827 ( .A(n12697), .B(n12891), .C(n2531), .Y(n6754) );
  NAND2X1 U4828 ( .A(ram[2317]), .B(n12891), .Y(n2531) );
  OAI21X1 U4829 ( .A(n12690), .B(n12891), .C(n2532), .Y(n6755) );
  NAND2X1 U4830 ( .A(ram[2318]), .B(n12891), .Y(n2532) );
  OAI21X1 U4831 ( .A(n12684), .B(n12891), .C(n2533), .Y(n6756) );
  NAND2X1 U4832 ( .A(ram[2319]), .B(n12891), .Y(n2533) );
  OAI21X1 U4834 ( .A(n12775), .B(n12890), .C(n2535), .Y(n6757) );
  NAND2X1 U4835 ( .A(ram[2320]), .B(n12890), .Y(n2535) );
  OAI21X1 U4836 ( .A(n12769), .B(n12890), .C(n2536), .Y(n6758) );
  NAND2X1 U4837 ( .A(ram[2321]), .B(n12890), .Y(n2536) );
  OAI21X1 U4838 ( .A(n12766), .B(n12890), .C(n2537), .Y(n6759) );
  NAND2X1 U4839 ( .A(ram[2322]), .B(n12890), .Y(n2537) );
  OAI21X1 U4840 ( .A(n12760), .B(n12890), .C(n2538), .Y(n6760) );
  NAND2X1 U4841 ( .A(ram[2323]), .B(n12890), .Y(n2538) );
  OAI21X1 U4842 ( .A(n12754), .B(n12890), .C(n2539), .Y(n6761) );
  NAND2X1 U4843 ( .A(ram[2324]), .B(n12890), .Y(n2539) );
  OAI21X1 U4844 ( .A(n12748), .B(n12890), .C(n2540), .Y(n6762) );
  NAND2X1 U4845 ( .A(ram[2325]), .B(n12890), .Y(n2540) );
  OAI21X1 U4846 ( .A(n12742), .B(n12890), .C(n2541), .Y(n6763) );
  NAND2X1 U4847 ( .A(ram[2326]), .B(n12890), .Y(n2541) );
  OAI21X1 U4848 ( .A(n12736), .B(n12890), .C(n2542), .Y(n6764) );
  NAND2X1 U4849 ( .A(ram[2327]), .B(n12890), .Y(n2542) );
  OAI21X1 U4850 ( .A(n12730), .B(n12890), .C(n2543), .Y(n6765) );
  NAND2X1 U4851 ( .A(ram[2328]), .B(n12890), .Y(n2543) );
  OAI21X1 U4852 ( .A(n12724), .B(n12890), .C(n2544), .Y(n6766) );
  NAND2X1 U4853 ( .A(ram[2329]), .B(n12890), .Y(n2544) );
  OAI21X1 U4854 ( .A(n12718), .B(n12890), .C(n2545), .Y(n6767) );
  NAND2X1 U4855 ( .A(ram[2330]), .B(n12890), .Y(n2545) );
  OAI21X1 U4856 ( .A(n12712), .B(n12890), .C(n2546), .Y(n6768) );
  NAND2X1 U4857 ( .A(ram[2331]), .B(n12890), .Y(n2546) );
  OAI21X1 U4858 ( .A(n12706), .B(n12890), .C(n2547), .Y(n6769) );
  NAND2X1 U4859 ( .A(ram[2332]), .B(n12890), .Y(n2547) );
  OAI21X1 U4860 ( .A(n12700), .B(n12890), .C(n2548), .Y(n6770) );
  NAND2X1 U4861 ( .A(ram[2333]), .B(n12890), .Y(n2548) );
  OAI21X1 U4862 ( .A(n12691), .B(n12890), .C(n2549), .Y(n6771) );
  NAND2X1 U4863 ( .A(ram[2334]), .B(n12890), .Y(n2549) );
  OAI21X1 U4864 ( .A(n12685), .B(n12890), .C(n2550), .Y(n6772) );
  NAND2X1 U4865 ( .A(ram[2335]), .B(n12890), .Y(n2550) );
  OAI21X1 U4867 ( .A(n12774), .B(n12889), .C(n2552), .Y(n6773) );
  NAND2X1 U4868 ( .A(ram[2336]), .B(n12889), .Y(n2552) );
  OAI21X1 U4869 ( .A(n12768), .B(n12889), .C(n2553), .Y(n6774) );
  NAND2X1 U4870 ( .A(ram[2337]), .B(n12889), .Y(n2553) );
  OAI21X1 U4871 ( .A(n12766), .B(n12889), .C(n2554), .Y(n6775) );
  NAND2X1 U4872 ( .A(ram[2338]), .B(n12889), .Y(n2554) );
  OAI21X1 U4873 ( .A(n12760), .B(n12889), .C(n2555), .Y(n6776) );
  NAND2X1 U4874 ( .A(ram[2339]), .B(n12889), .Y(n2555) );
  OAI21X1 U4875 ( .A(n12754), .B(n12889), .C(n2556), .Y(n6777) );
  NAND2X1 U4876 ( .A(ram[2340]), .B(n12889), .Y(n2556) );
  OAI21X1 U4877 ( .A(n12748), .B(n12889), .C(n2557), .Y(n6778) );
  NAND2X1 U4878 ( .A(ram[2341]), .B(n12889), .Y(n2557) );
  OAI21X1 U4879 ( .A(n12742), .B(n12889), .C(n2558), .Y(n6779) );
  NAND2X1 U4880 ( .A(ram[2342]), .B(n12889), .Y(n2558) );
  OAI21X1 U4881 ( .A(n12736), .B(n12889), .C(n2559), .Y(n6780) );
  NAND2X1 U4882 ( .A(ram[2343]), .B(n12889), .Y(n2559) );
  OAI21X1 U4883 ( .A(n12730), .B(n12889), .C(n2560), .Y(n6781) );
  NAND2X1 U4884 ( .A(ram[2344]), .B(n12889), .Y(n2560) );
  OAI21X1 U4885 ( .A(n12724), .B(n12889), .C(n2561), .Y(n6782) );
  NAND2X1 U4886 ( .A(ram[2345]), .B(n12889), .Y(n2561) );
  OAI21X1 U4887 ( .A(n12718), .B(n12889), .C(n2562), .Y(n6783) );
  NAND2X1 U4888 ( .A(ram[2346]), .B(n12889), .Y(n2562) );
  OAI21X1 U4889 ( .A(n12712), .B(n12889), .C(n2563), .Y(n6784) );
  NAND2X1 U4890 ( .A(ram[2347]), .B(n12889), .Y(n2563) );
  OAI21X1 U4891 ( .A(n12706), .B(n12889), .C(n2564), .Y(n6785) );
  NAND2X1 U4892 ( .A(ram[2348]), .B(n12889), .Y(n2564) );
  OAI21X1 U4893 ( .A(n12700), .B(n12889), .C(n2565), .Y(n6786) );
  NAND2X1 U4894 ( .A(ram[2349]), .B(n12889), .Y(n2565) );
  OAI21X1 U4895 ( .A(n12690), .B(n12889), .C(n2566), .Y(n6787) );
  NAND2X1 U4896 ( .A(ram[2350]), .B(n12889), .Y(n2566) );
  OAI21X1 U4897 ( .A(n12684), .B(n12889), .C(n2567), .Y(n6788) );
  NAND2X1 U4898 ( .A(ram[2351]), .B(n12889), .Y(n2567) );
  OAI21X1 U4900 ( .A(n12779), .B(n12888), .C(n2569), .Y(n6789) );
  NAND2X1 U4901 ( .A(ram[2352]), .B(n12888), .Y(n2569) );
  OAI21X1 U4902 ( .A(n12773), .B(n12888), .C(n2570), .Y(n6790) );
  NAND2X1 U4903 ( .A(ram[2353]), .B(n12888), .Y(n2570) );
  OAI21X1 U4904 ( .A(n12766), .B(n12888), .C(n2571), .Y(n6791) );
  NAND2X1 U4905 ( .A(ram[2354]), .B(n12888), .Y(n2571) );
  OAI21X1 U4906 ( .A(n12760), .B(n12888), .C(n2572), .Y(n6792) );
  NAND2X1 U4907 ( .A(ram[2355]), .B(n12888), .Y(n2572) );
  OAI21X1 U4908 ( .A(n12754), .B(n12888), .C(n2573), .Y(n6793) );
  NAND2X1 U4909 ( .A(ram[2356]), .B(n12888), .Y(n2573) );
  OAI21X1 U4910 ( .A(n12748), .B(n12888), .C(n2574), .Y(n6794) );
  NAND2X1 U4911 ( .A(ram[2357]), .B(n12888), .Y(n2574) );
  OAI21X1 U4912 ( .A(n12742), .B(n12888), .C(n2575), .Y(n6795) );
  NAND2X1 U4913 ( .A(ram[2358]), .B(n12888), .Y(n2575) );
  OAI21X1 U4914 ( .A(n12736), .B(n12888), .C(n2576), .Y(n6796) );
  NAND2X1 U4915 ( .A(ram[2359]), .B(n12888), .Y(n2576) );
  OAI21X1 U4916 ( .A(n12730), .B(n12888), .C(n2577), .Y(n6797) );
  NAND2X1 U4917 ( .A(ram[2360]), .B(n12888), .Y(n2577) );
  OAI21X1 U4918 ( .A(n12724), .B(n12888), .C(n2578), .Y(n6798) );
  NAND2X1 U4919 ( .A(ram[2361]), .B(n12888), .Y(n2578) );
  OAI21X1 U4920 ( .A(n12718), .B(n12888), .C(n2579), .Y(n6799) );
  NAND2X1 U4921 ( .A(ram[2362]), .B(n12888), .Y(n2579) );
  OAI21X1 U4922 ( .A(n12712), .B(n12888), .C(n2580), .Y(n6800) );
  NAND2X1 U4923 ( .A(ram[2363]), .B(n12888), .Y(n2580) );
  OAI21X1 U4924 ( .A(n12706), .B(n12888), .C(n2581), .Y(n6801) );
  NAND2X1 U4925 ( .A(ram[2364]), .B(n12888), .Y(n2581) );
  OAI21X1 U4926 ( .A(n12700), .B(n12888), .C(n2582), .Y(n6802) );
  NAND2X1 U4927 ( .A(ram[2365]), .B(n12888), .Y(n2582) );
  OAI21X1 U4928 ( .A(n12695), .B(n12888), .C(n2583), .Y(n6803) );
  NAND2X1 U4929 ( .A(ram[2366]), .B(n12888), .Y(n2583) );
  OAI21X1 U4930 ( .A(n12689), .B(n12888), .C(n2584), .Y(n6804) );
  NAND2X1 U4931 ( .A(ram[2367]), .B(n12888), .Y(n2584) );
  OAI21X1 U4933 ( .A(n12778), .B(n12887), .C(n2586), .Y(n6805) );
  NAND2X1 U4934 ( .A(ram[2368]), .B(n12887), .Y(n2586) );
  OAI21X1 U4935 ( .A(n12772), .B(n12887), .C(n2587), .Y(n6806) );
  NAND2X1 U4936 ( .A(ram[2369]), .B(n12887), .Y(n2587) );
  OAI21X1 U4937 ( .A(n12764), .B(n12887), .C(n2588), .Y(n6807) );
  NAND2X1 U4938 ( .A(ram[2370]), .B(n12887), .Y(n2588) );
  OAI21X1 U4939 ( .A(n12758), .B(n12887), .C(n2589), .Y(n6808) );
  NAND2X1 U4940 ( .A(ram[2371]), .B(n12887), .Y(n2589) );
  OAI21X1 U4941 ( .A(n12752), .B(n12887), .C(n2590), .Y(n6809) );
  NAND2X1 U4942 ( .A(ram[2372]), .B(n12887), .Y(n2590) );
  OAI21X1 U4943 ( .A(n12746), .B(n12887), .C(n2591), .Y(n6810) );
  NAND2X1 U4944 ( .A(ram[2373]), .B(n12887), .Y(n2591) );
  OAI21X1 U4945 ( .A(n12740), .B(n12887), .C(n2592), .Y(n6811) );
  NAND2X1 U4946 ( .A(ram[2374]), .B(n12887), .Y(n2592) );
  OAI21X1 U4947 ( .A(n12734), .B(n12887), .C(n2593), .Y(n6812) );
  NAND2X1 U4948 ( .A(ram[2375]), .B(n12887), .Y(n2593) );
  OAI21X1 U4949 ( .A(n12728), .B(n12887), .C(n2594), .Y(n6813) );
  NAND2X1 U4950 ( .A(ram[2376]), .B(n12887), .Y(n2594) );
  OAI21X1 U4951 ( .A(n12722), .B(n12887), .C(n2595), .Y(n6814) );
  NAND2X1 U4952 ( .A(ram[2377]), .B(n12887), .Y(n2595) );
  OAI21X1 U4953 ( .A(n12716), .B(n12887), .C(n2596), .Y(n6815) );
  NAND2X1 U4954 ( .A(ram[2378]), .B(n12887), .Y(n2596) );
  OAI21X1 U4955 ( .A(n12710), .B(n12887), .C(n2597), .Y(n6816) );
  NAND2X1 U4956 ( .A(ram[2379]), .B(n12887), .Y(n2597) );
  OAI21X1 U4957 ( .A(n12704), .B(n12887), .C(n2598), .Y(n6817) );
  NAND2X1 U4958 ( .A(ram[2380]), .B(n12887), .Y(n2598) );
  OAI21X1 U4959 ( .A(n12698), .B(n12887), .C(n2599), .Y(n6818) );
  NAND2X1 U4960 ( .A(ram[2381]), .B(n12887), .Y(n2599) );
  OAI21X1 U4961 ( .A(n12694), .B(n12887), .C(n2600), .Y(n6819) );
  NAND2X1 U4962 ( .A(ram[2382]), .B(n12887), .Y(n2600) );
  OAI21X1 U4963 ( .A(n12688), .B(n12887), .C(n2601), .Y(n6820) );
  NAND2X1 U4964 ( .A(ram[2383]), .B(n12887), .Y(n2601) );
  OAI21X1 U4966 ( .A(n12777), .B(n12886), .C(n2603), .Y(n6821) );
  NAND2X1 U4967 ( .A(ram[2384]), .B(n12886), .Y(n2603) );
  OAI21X1 U4968 ( .A(n12771), .B(n12886), .C(n2604), .Y(n6822) );
  NAND2X1 U4969 ( .A(ram[2385]), .B(n12886), .Y(n2604) );
  OAI21X1 U4970 ( .A(n12762), .B(n12886), .C(n2605), .Y(n6823) );
  NAND2X1 U4971 ( .A(ram[2386]), .B(n12886), .Y(n2605) );
  OAI21X1 U4972 ( .A(n12756), .B(n12886), .C(n2606), .Y(n6824) );
  NAND2X1 U4973 ( .A(ram[2387]), .B(n12886), .Y(n2606) );
  OAI21X1 U4974 ( .A(n12750), .B(n12886), .C(n2607), .Y(n6825) );
  NAND2X1 U4975 ( .A(ram[2388]), .B(n12886), .Y(n2607) );
  OAI21X1 U4976 ( .A(n12744), .B(n12886), .C(n2608), .Y(n6826) );
  NAND2X1 U4977 ( .A(ram[2389]), .B(n12886), .Y(n2608) );
  OAI21X1 U4978 ( .A(n12738), .B(n12886), .C(n2609), .Y(n6827) );
  NAND2X1 U4979 ( .A(ram[2390]), .B(n12886), .Y(n2609) );
  OAI21X1 U4980 ( .A(n12732), .B(n12886), .C(n2610), .Y(n6828) );
  NAND2X1 U4981 ( .A(ram[2391]), .B(n12886), .Y(n2610) );
  OAI21X1 U4982 ( .A(n12726), .B(n12886), .C(n2611), .Y(n6829) );
  NAND2X1 U4983 ( .A(ram[2392]), .B(n12886), .Y(n2611) );
  OAI21X1 U4984 ( .A(n12720), .B(n12886), .C(n2612), .Y(n6830) );
  NAND2X1 U4985 ( .A(ram[2393]), .B(n12886), .Y(n2612) );
  OAI21X1 U4986 ( .A(n12714), .B(n12886), .C(n2613), .Y(n6831) );
  NAND2X1 U4987 ( .A(ram[2394]), .B(n12886), .Y(n2613) );
  OAI21X1 U4988 ( .A(n12708), .B(n12886), .C(n2614), .Y(n6832) );
  NAND2X1 U4989 ( .A(ram[2395]), .B(n12886), .Y(n2614) );
  OAI21X1 U4990 ( .A(n12702), .B(n12886), .C(n2615), .Y(n6833) );
  NAND2X1 U4991 ( .A(ram[2396]), .B(n12886), .Y(n2615) );
  OAI21X1 U4992 ( .A(n12696), .B(n12886), .C(n2616), .Y(n6834) );
  NAND2X1 U4993 ( .A(ram[2397]), .B(n12886), .Y(n2616) );
  OAI21X1 U4994 ( .A(n12693), .B(n12886), .C(n2617), .Y(n6835) );
  NAND2X1 U4995 ( .A(ram[2398]), .B(n12886), .Y(n2617) );
  OAI21X1 U4996 ( .A(n12687), .B(n12886), .C(n2618), .Y(n6836) );
  NAND2X1 U4997 ( .A(ram[2399]), .B(n12886), .Y(n2618) );
  OAI21X1 U4999 ( .A(n12774), .B(n12885), .C(n2620), .Y(n6837) );
  NAND2X1 U5000 ( .A(ram[2400]), .B(n12885), .Y(n2620) );
  OAI21X1 U5001 ( .A(n12768), .B(n12885), .C(n2621), .Y(n6838) );
  NAND2X1 U5002 ( .A(ram[2401]), .B(n12885), .Y(n2621) );
  OAI21X1 U5003 ( .A(n12763), .B(n12885), .C(n2622), .Y(n6839) );
  NAND2X1 U5004 ( .A(ram[2402]), .B(n12885), .Y(n2622) );
  OAI21X1 U5005 ( .A(n12757), .B(n12885), .C(n2623), .Y(n6840) );
  NAND2X1 U5006 ( .A(ram[2403]), .B(n12885), .Y(n2623) );
  OAI21X1 U5007 ( .A(n12751), .B(n12885), .C(n2624), .Y(n6841) );
  NAND2X1 U5008 ( .A(ram[2404]), .B(n12885), .Y(n2624) );
  OAI21X1 U5009 ( .A(n12745), .B(n12885), .C(n2625), .Y(n6842) );
  NAND2X1 U5010 ( .A(ram[2405]), .B(n12885), .Y(n2625) );
  OAI21X1 U5011 ( .A(n12739), .B(n12885), .C(n2626), .Y(n6843) );
  NAND2X1 U5012 ( .A(ram[2406]), .B(n12885), .Y(n2626) );
  OAI21X1 U5013 ( .A(n12733), .B(n12885), .C(n2627), .Y(n6844) );
  NAND2X1 U5014 ( .A(ram[2407]), .B(n12885), .Y(n2627) );
  OAI21X1 U5015 ( .A(n12727), .B(n12885), .C(n2628), .Y(n6845) );
  NAND2X1 U5016 ( .A(ram[2408]), .B(n12885), .Y(n2628) );
  OAI21X1 U5017 ( .A(n12721), .B(n12885), .C(n2629), .Y(n6846) );
  NAND2X1 U5018 ( .A(ram[2409]), .B(n12885), .Y(n2629) );
  OAI21X1 U5019 ( .A(n12715), .B(n12885), .C(n2630), .Y(n6847) );
  NAND2X1 U5020 ( .A(ram[2410]), .B(n12885), .Y(n2630) );
  OAI21X1 U5021 ( .A(n12709), .B(n12885), .C(n2631), .Y(n6848) );
  NAND2X1 U5022 ( .A(ram[2411]), .B(n12885), .Y(n2631) );
  OAI21X1 U5023 ( .A(n12703), .B(n12885), .C(n2632), .Y(n6849) );
  NAND2X1 U5024 ( .A(ram[2412]), .B(n12885), .Y(n2632) );
  OAI21X1 U5025 ( .A(n12697), .B(n12885), .C(n2633), .Y(n6850) );
  NAND2X1 U5026 ( .A(ram[2413]), .B(n12885), .Y(n2633) );
  OAI21X1 U5027 ( .A(n12690), .B(n12885), .C(n2634), .Y(n6851) );
  NAND2X1 U5028 ( .A(ram[2414]), .B(n12885), .Y(n2634) );
  OAI21X1 U5029 ( .A(n12684), .B(n12885), .C(n2635), .Y(n6852) );
  NAND2X1 U5030 ( .A(ram[2415]), .B(n12885), .Y(n2635) );
  OAI21X1 U5032 ( .A(n12776), .B(n12884), .C(n2637), .Y(n6853) );
  NAND2X1 U5033 ( .A(ram[2416]), .B(n12884), .Y(n2637) );
  OAI21X1 U5034 ( .A(n12770), .B(n12884), .C(n2638), .Y(n6854) );
  NAND2X1 U5035 ( .A(ram[2417]), .B(n12884), .Y(n2638) );
  OAI21X1 U5036 ( .A(n12762), .B(n12884), .C(n2639), .Y(n6855) );
  NAND2X1 U5037 ( .A(ram[2418]), .B(n12884), .Y(n2639) );
  OAI21X1 U5038 ( .A(n12756), .B(n12884), .C(n2640), .Y(n6856) );
  NAND2X1 U5039 ( .A(ram[2419]), .B(n12884), .Y(n2640) );
  OAI21X1 U5040 ( .A(n12750), .B(n12884), .C(n2641), .Y(n6857) );
  NAND2X1 U5041 ( .A(ram[2420]), .B(n12884), .Y(n2641) );
  OAI21X1 U5042 ( .A(n12744), .B(n12884), .C(n2642), .Y(n6858) );
  NAND2X1 U5043 ( .A(ram[2421]), .B(n12884), .Y(n2642) );
  OAI21X1 U5044 ( .A(n12738), .B(n12884), .C(n2643), .Y(n6859) );
  NAND2X1 U5045 ( .A(ram[2422]), .B(n12884), .Y(n2643) );
  OAI21X1 U5046 ( .A(n12732), .B(n12884), .C(n2644), .Y(n6860) );
  NAND2X1 U5047 ( .A(ram[2423]), .B(n12884), .Y(n2644) );
  OAI21X1 U5048 ( .A(n12726), .B(n12884), .C(n2645), .Y(n6861) );
  NAND2X1 U5049 ( .A(ram[2424]), .B(n12884), .Y(n2645) );
  OAI21X1 U5050 ( .A(n12720), .B(n12884), .C(n2646), .Y(n6862) );
  NAND2X1 U5051 ( .A(ram[2425]), .B(n12884), .Y(n2646) );
  OAI21X1 U5052 ( .A(n12714), .B(n12884), .C(n2647), .Y(n6863) );
  NAND2X1 U5053 ( .A(ram[2426]), .B(n12884), .Y(n2647) );
  OAI21X1 U5054 ( .A(n12708), .B(n12884), .C(n2648), .Y(n6864) );
  NAND2X1 U5055 ( .A(ram[2427]), .B(n12884), .Y(n2648) );
  OAI21X1 U5056 ( .A(n12702), .B(n12884), .C(n2649), .Y(n6865) );
  NAND2X1 U5057 ( .A(ram[2428]), .B(n12884), .Y(n2649) );
  OAI21X1 U5058 ( .A(n12696), .B(n12884), .C(n2650), .Y(n6866) );
  NAND2X1 U5059 ( .A(ram[2429]), .B(n12884), .Y(n2650) );
  OAI21X1 U5060 ( .A(n12692), .B(n12884), .C(n2651), .Y(n6867) );
  NAND2X1 U5061 ( .A(ram[2430]), .B(n12884), .Y(n2651) );
  OAI21X1 U5062 ( .A(n12686), .B(n12884), .C(n2652), .Y(n6868) );
  NAND2X1 U5063 ( .A(ram[2431]), .B(n12884), .Y(n2652) );
  OAI21X1 U5065 ( .A(n12775), .B(n12883), .C(n2654), .Y(n6869) );
  NAND2X1 U5066 ( .A(ram[2432]), .B(n12883), .Y(n2654) );
  OAI21X1 U5067 ( .A(n12769), .B(n12883), .C(n2655), .Y(n6870) );
  NAND2X1 U5068 ( .A(ram[2433]), .B(n12883), .Y(n2655) );
  OAI21X1 U5069 ( .A(n12763), .B(n12883), .C(n2656), .Y(n6871) );
  NAND2X1 U5070 ( .A(ram[2434]), .B(n12883), .Y(n2656) );
  OAI21X1 U5071 ( .A(n12757), .B(n12883), .C(n2657), .Y(n6872) );
  NAND2X1 U5072 ( .A(ram[2435]), .B(n12883), .Y(n2657) );
  OAI21X1 U5073 ( .A(n12751), .B(n12883), .C(n2658), .Y(n6873) );
  NAND2X1 U5074 ( .A(ram[2436]), .B(n12883), .Y(n2658) );
  OAI21X1 U5075 ( .A(n12745), .B(n12883), .C(n2659), .Y(n6874) );
  NAND2X1 U5076 ( .A(ram[2437]), .B(n12883), .Y(n2659) );
  OAI21X1 U5077 ( .A(n12739), .B(n12883), .C(n2660), .Y(n6875) );
  NAND2X1 U5078 ( .A(ram[2438]), .B(n12883), .Y(n2660) );
  OAI21X1 U5079 ( .A(n12733), .B(n12883), .C(n2661), .Y(n6876) );
  NAND2X1 U5080 ( .A(ram[2439]), .B(n12883), .Y(n2661) );
  OAI21X1 U5081 ( .A(n12727), .B(n12883), .C(n2662), .Y(n6877) );
  NAND2X1 U5082 ( .A(ram[2440]), .B(n12883), .Y(n2662) );
  OAI21X1 U5083 ( .A(n12721), .B(n12883), .C(n2663), .Y(n6878) );
  NAND2X1 U5084 ( .A(ram[2441]), .B(n12883), .Y(n2663) );
  OAI21X1 U5085 ( .A(n12715), .B(n12883), .C(n2664), .Y(n6879) );
  NAND2X1 U5086 ( .A(ram[2442]), .B(n12883), .Y(n2664) );
  OAI21X1 U5087 ( .A(n12709), .B(n12883), .C(n2665), .Y(n6880) );
  NAND2X1 U5088 ( .A(ram[2443]), .B(n12883), .Y(n2665) );
  OAI21X1 U5089 ( .A(n12703), .B(n12883), .C(n2666), .Y(n6881) );
  NAND2X1 U5090 ( .A(ram[2444]), .B(n12883), .Y(n2666) );
  OAI21X1 U5091 ( .A(n12697), .B(n12883), .C(n2667), .Y(n6882) );
  NAND2X1 U5092 ( .A(ram[2445]), .B(n12883), .Y(n2667) );
  OAI21X1 U5093 ( .A(n12691), .B(n12883), .C(n2668), .Y(n6883) );
  NAND2X1 U5094 ( .A(ram[2446]), .B(n12883), .Y(n2668) );
  OAI21X1 U5095 ( .A(n12685), .B(n12883), .C(n2669), .Y(n6884) );
  NAND2X1 U5096 ( .A(ram[2447]), .B(n12883), .Y(n2669) );
  OAI21X1 U5098 ( .A(n12774), .B(n12882), .C(n2671), .Y(n6885) );
  NAND2X1 U5099 ( .A(ram[2448]), .B(n12882), .Y(n2671) );
  OAI21X1 U5100 ( .A(n12768), .B(n12882), .C(n2672), .Y(n6886) );
  NAND2X1 U5101 ( .A(ram[2449]), .B(n12882), .Y(n2672) );
  OAI21X1 U5102 ( .A(n12767), .B(n12882), .C(n2673), .Y(n6887) );
  NAND2X1 U5103 ( .A(ram[2450]), .B(n12882), .Y(n2673) );
  OAI21X1 U5104 ( .A(n12761), .B(n12882), .C(n2674), .Y(n6888) );
  NAND2X1 U5105 ( .A(ram[2451]), .B(n12882), .Y(n2674) );
  OAI21X1 U5106 ( .A(n12755), .B(n12882), .C(n2675), .Y(n6889) );
  NAND2X1 U5107 ( .A(ram[2452]), .B(n12882), .Y(n2675) );
  OAI21X1 U5108 ( .A(n12749), .B(n12882), .C(n2676), .Y(n6890) );
  NAND2X1 U5109 ( .A(ram[2453]), .B(n12882), .Y(n2676) );
  OAI21X1 U5110 ( .A(n12743), .B(n12882), .C(n2677), .Y(n6891) );
  NAND2X1 U5111 ( .A(ram[2454]), .B(n12882), .Y(n2677) );
  OAI21X1 U5112 ( .A(n12737), .B(n12882), .C(n2678), .Y(n6892) );
  NAND2X1 U5113 ( .A(ram[2455]), .B(n12882), .Y(n2678) );
  OAI21X1 U5114 ( .A(n12731), .B(n12882), .C(n2679), .Y(n6893) );
  NAND2X1 U5115 ( .A(ram[2456]), .B(n12882), .Y(n2679) );
  OAI21X1 U5116 ( .A(n12725), .B(n12882), .C(n2680), .Y(n6894) );
  NAND2X1 U5117 ( .A(ram[2457]), .B(n12882), .Y(n2680) );
  OAI21X1 U5118 ( .A(n12719), .B(n12882), .C(n2681), .Y(n6895) );
  NAND2X1 U5119 ( .A(ram[2458]), .B(n12882), .Y(n2681) );
  OAI21X1 U5120 ( .A(n12713), .B(n12882), .C(n2682), .Y(n6896) );
  NAND2X1 U5121 ( .A(ram[2459]), .B(n12882), .Y(n2682) );
  OAI21X1 U5122 ( .A(n12707), .B(n12882), .C(n2683), .Y(n6897) );
  NAND2X1 U5123 ( .A(ram[2460]), .B(n12882), .Y(n2683) );
  OAI21X1 U5124 ( .A(n12701), .B(n12882), .C(n2684), .Y(n6898) );
  NAND2X1 U5125 ( .A(ram[2461]), .B(n12882), .Y(n2684) );
  OAI21X1 U5126 ( .A(n12690), .B(n12882), .C(n2685), .Y(n6899) );
  NAND2X1 U5127 ( .A(ram[2462]), .B(n12882), .Y(n2685) );
  OAI21X1 U5128 ( .A(n12684), .B(n12882), .C(n2686), .Y(n6900) );
  NAND2X1 U5129 ( .A(ram[2463]), .B(n12882), .Y(n2686) );
  OAI21X1 U5131 ( .A(n12774), .B(n12881), .C(n2688), .Y(n6901) );
  NAND2X1 U5132 ( .A(ram[2464]), .B(n12881), .Y(n2688) );
  OAI21X1 U5133 ( .A(n12768), .B(n12881), .C(n2689), .Y(n6902) );
  NAND2X1 U5134 ( .A(ram[2465]), .B(n12881), .Y(n2689) );
  OAI21X1 U5135 ( .A(n12766), .B(n12881), .C(n2690), .Y(n6903) );
  NAND2X1 U5136 ( .A(ram[2466]), .B(n12881), .Y(n2690) );
  OAI21X1 U5137 ( .A(n12760), .B(n12881), .C(n2691), .Y(n6904) );
  NAND2X1 U5138 ( .A(ram[2467]), .B(n12881), .Y(n2691) );
  OAI21X1 U5139 ( .A(n12754), .B(n12881), .C(n2692), .Y(n6905) );
  NAND2X1 U5140 ( .A(ram[2468]), .B(n12881), .Y(n2692) );
  OAI21X1 U5141 ( .A(n12748), .B(n12881), .C(n2693), .Y(n6906) );
  NAND2X1 U5142 ( .A(ram[2469]), .B(n12881), .Y(n2693) );
  OAI21X1 U5143 ( .A(n12742), .B(n12881), .C(n2694), .Y(n6907) );
  NAND2X1 U5144 ( .A(ram[2470]), .B(n12881), .Y(n2694) );
  OAI21X1 U5145 ( .A(n12736), .B(n12881), .C(n2695), .Y(n6908) );
  NAND2X1 U5146 ( .A(ram[2471]), .B(n12881), .Y(n2695) );
  OAI21X1 U5147 ( .A(n12730), .B(n12881), .C(n2696), .Y(n6909) );
  NAND2X1 U5148 ( .A(ram[2472]), .B(n12881), .Y(n2696) );
  OAI21X1 U5149 ( .A(n12724), .B(n12881), .C(n2697), .Y(n6910) );
  NAND2X1 U5150 ( .A(ram[2473]), .B(n12881), .Y(n2697) );
  OAI21X1 U5151 ( .A(n12718), .B(n12881), .C(n2698), .Y(n6911) );
  NAND2X1 U5152 ( .A(ram[2474]), .B(n12881), .Y(n2698) );
  OAI21X1 U5153 ( .A(n12712), .B(n12881), .C(n2699), .Y(n6912) );
  NAND2X1 U5154 ( .A(ram[2475]), .B(n12881), .Y(n2699) );
  OAI21X1 U5155 ( .A(n12706), .B(n12881), .C(n2700), .Y(n6913) );
  NAND2X1 U5156 ( .A(ram[2476]), .B(n12881), .Y(n2700) );
  OAI21X1 U5157 ( .A(n12700), .B(n12881), .C(n2701), .Y(n6914) );
  NAND2X1 U5158 ( .A(ram[2477]), .B(n12881), .Y(n2701) );
  OAI21X1 U5159 ( .A(n12690), .B(n12881), .C(n2702), .Y(n6915) );
  NAND2X1 U5160 ( .A(ram[2478]), .B(n12881), .Y(n2702) );
  OAI21X1 U5161 ( .A(n12684), .B(n12881), .C(n2703), .Y(n6916) );
  NAND2X1 U5162 ( .A(ram[2479]), .B(n12881), .Y(n2703) );
  OAI21X1 U5164 ( .A(n12776), .B(n12880), .C(n2705), .Y(n6917) );
  NAND2X1 U5165 ( .A(ram[2480]), .B(n12880), .Y(n2705) );
  OAI21X1 U5166 ( .A(n12770), .B(n12880), .C(n2706), .Y(n6918) );
  NAND2X1 U5167 ( .A(ram[2481]), .B(n12880), .Y(n2706) );
  OAI21X1 U5168 ( .A(n12762), .B(n12880), .C(n2707), .Y(n6919) );
  NAND2X1 U5169 ( .A(ram[2482]), .B(n12880), .Y(n2707) );
  OAI21X1 U5170 ( .A(n12756), .B(n12880), .C(n2708), .Y(n6920) );
  NAND2X1 U5171 ( .A(ram[2483]), .B(n12880), .Y(n2708) );
  OAI21X1 U5172 ( .A(n12750), .B(n12880), .C(n2709), .Y(n6921) );
  NAND2X1 U5173 ( .A(ram[2484]), .B(n12880), .Y(n2709) );
  OAI21X1 U5174 ( .A(n12744), .B(n12880), .C(n2710), .Y(n6922) );
  NAND2X1 U5175 ( .A(ram[2485]), .B(n12880), .Y(n2710) );
  OAI21X1 U5176 ( .A(n12738), .B(n12880), .C(n2711), .Y(n6923) );
  NAND2X1 U5177 ( .A(ram[2486]), .B(n12880), .Y(n2711) );
  OAI21X1 U5178 ( .A(n12732), .B(n12880), .C(n2712), .Y(n6924) );
  NAND2X1 U5179 ( .A(ram[2487]), .B(n12880), .Y(n2712) );
  OAI21X1 U5180 ( .A(n12726), .B(n12880), .C(n2713), .Y(n6925) );
  NAND2X1 U5181 ( .A(ram[2488]), .B(n12880), .Y(n2713) );
  OAI21X1 U5182 ( .A(n12720), .B(n12880), .C(n2714), .Y(n6926) );
  NAND2X1 U5183 ( .A(ram[2489]), .B(n12880), .Y(n2714) );
  OAI21X1 U5184 ( .A(n12714), .B(n12880), .C(n2715), .Y(n6927) );
  NAND2X1 U5185 ( .A(ram[2490]), .B(n12880), .Y(n2715) );
  OAI21X1 U5186 ( .A(n12708), .B(n12880), .C(n2716), .Y(n6928) );
  NAND2X1 U5187 ( .A(ram[2491]), .B(n12880), .Y(n2716) );
  OAI21X1 U5188 ( .A(n12702), .B(n12880), .C(n2717), .Y(n6929) );
  NAND2X1 U5189 ( .A(ram[2492]), .B(n12880), .Y(n2717) );
  OAI21X1 U5190 ( .A(n12696), .B(n12880), .C(n2718), .Y(n6930) );
  NAND2X1 U5191 ( .A(ram[2493]), .B(n12880), .Y(n2718) );
  OAI21X1 U5192 ( .A(n12692), .B(n12880), .C(n2719), .Y(n6931) );
  NAND2X1 U5193 ( .A(ram[2494]), .B(n12880), .Y(n2719) );
  OAI21X1 U5194 ( .A(n12686), .B(n12880), .C(n2720), .Y(n6932) );
  NAND2X1 U5195 ( .A(ram[2495]), .B(n12880), .Y(n2720) );
  OAI21X1 U5197 ( .A(n12775), .B(n12879), .C(n2722), .Y(n6933) );
  NAND2X1 U5198 ( .A(ram[2496]), .B(n12879), .Y(n2722) );
  OAI21X1 U5199 ( .A(n12769), .B(n12879), .C(n2723), .Y(n6934) );
  NAND2X1 U5200 ( .A(ram[2497]), .B(n12879), .Y(n2723) );
  OAI21X1 U5201 ( .A(n12766), .B(n12879), .C(n2724), .Y(n6935) );
  NAND2X1 U5202 ( .A(ram[2498]), .B(n12879), .Y(n2724) );
  OAI21X1 U5203 ( .A(n12760), .B(n12879), .C(n2725), .Y(n6936) );
  NAND2X1 U5204 ( .A(ram[2499]), .B(n12879), .Y(n2725) );
  OAI21X1 U5205 ( .A(n12754), .B(n12879), .C(n2726), .Y(n6937) );
  NAND2X1 U5206 ( .A(ram[2500]), .B(n12879), .Y(n2726) );
  OAI21X1 U5207 ( .A(n12748), .B(n12879), .C(n2727), .Y(n6938) );
  NAND2X1 U5208 ( .A(ram[2501]), .B(n12879), .Y(n2727) );
  OAI21X1 U5209 ( .A(n12742), .B(n12879), .C(n2728), .Y(n6939) );
  NAND2X1 U5210 ( .A(ram[2502]), .B(n12879), .Y(n2728) );
  OAI21X1 U5211 ( .A(n12736), .B(n12879), .C(n2729), .Y(n6940) );
  NAND2X1 U5212 ( .A(ram[2503]), .B(n12879), .Y(n2729) );
  OAI21X1 U5213 ( .A(n12730), .B(n12879), .C(n2730), .Y(n6941) );
  NAND2X1 U5214 ( .A(ram[2504]), .B(n12879), .Y(n2730) );
  OAI21X1 U5215 ( .A(n12724), .B(n12879), .C(n2731), .Y(n6942) );
  NAND2X1 U5216 ( .A(ram[2505]), .B(n12879), .Y(n2731) );
  OAI21X1 U5217 ( .A(n12718), .B(n12879), .C(n2732), .Y(n6943) );
  NAND2X1 U5218 ( .A(ram[2506]), .B(n12879), .Y(n2732) );
  OAI21X1 U5219 ( .A(n12712), .B(n12879), .C(n2733), .Y(n6944) );
  NAND2X1 U5220 ( .A(ram[2507]), .B(n12879), .Y(n2733) );
  OAI21X1 U5221 ( .A(n12706), .B(n12879), .C(n2734), .Y(n6945) );
  NAND2X1 U5222 ( .A(ram[2508]), .B(n12879), .Y(n2734) );
  OAI21X1 U5223 ( .A(n12700), .B(n12879), .C(n2735), .Y(n6946) );
  NAND2X1 U5224 ( .A(ram[2509]), .B(n12879), .Y(n2735) );
  OAI21X1 U5225 ( .A(n12691), .B(n12879), .C(n2736), .Y(n6947) );
  NAND2X1 U5226 ( .A(ram[2510]), .B(n12879), .Y(n2736) );
  OAI21X1 U5227 ( .A(n12685), .B(n12879), .C(n2737), .Y(n6948) );
  NAND2X1 U5228 ( .A(ram[2511]), .B(n12879), .Y(n2737) );
  OAI21X1 U5230 ( .A(n12775), .B(n12878), .C(n2739), .Y(n6949) );
  NAND2X1 U5231 ( .A(ram[2512]), .B(n12878), .Y(n2739) );
  OAI21X1 U5232 ( .A(n12769), .B(n12878), .C(n2740), .Y(n6950) );
  NAND2X1 U5233 ( .A(ram[2513]), .B(n12878), .Y(n2740) );
  OAI21X1 U5234 ( .A(n12762), .B(n12878), .C(n2741), .Y(n6951) );
  NAND2X1 U5235 ( .A(ram[2514]), .B(n12878), .Y(n2741) );
  OAI21X1 U5236 ( .A(n12756), .B(n12878), .C(n2742), .Y(n6952) );
  NAND2X1 U5237 ( .A(ram[2515]), .B(n12878), .Y(n2742) );
  OAI21X1 U5238 ( .A(n12750), .B(n12878), .C(n2743), .Y(n6953) );
  NAND2X1 U5239 ( .A(ram[2516]), .B(n12878), .Y(n2743) );
  OAI21X1 U5240 ( .A(n12744), .B(n12878), .C(n2744), .Y(n6954) );
  NAND2X1 U5241 ( .A(ram[2517]), .B(n12878), .Y(n2744) );
  OAI21X1 U5242 ( .A(n12738), .B(n12878), .C(n2745), .Y(n6955) );
  NAND2X1 U5243 ( .A(ram[2518]), .B(n12878), .Y(n2745) );
  OAI21X1 U5244 ( .A(n12732), .B(n12878), .C(n2746), .Y(n6956) );
  NAND2X1 U5245 ( .A(ram[2519]), .B(n12878), .Y(n2746) );
  OAI21X1 U5246 ( .A(n12726), .B(n12878), .C(n2747), .Y(n6957) );
  NAND2X1 U5247 ( .A(ram[2520]), .B(n12878), .Y(n2747) );
  OAI21X1 U5248 ( .A(n12720), .B(n12878), .C(n2748), .Y(n6958) );
  NAND2X1 U5249 ( .A(ram[2521]), .B(n12878), .Y(n2748) );
  OAI21X1 U5250 ( .A(n12714), .B(n12878), .C(n2749), .Y(n6959) );
  NAND2X1 U5251 ( .A(ram[2522]), .B(n12878), .Y(n2749) );
  OAI21X1 U5252 ( .A(n12708), .B(n12878), .C(n2750), .Y(n6960) );
  NAND2X1 U5253 ( .A(ram[2523]), .B(n12878), .Y(n2750) );
  OAI21X1 U5254 ( .A(n12702), .B(n12878), .C(n2751), .Y(n6961) );
  NAND2X1 U5255 ( .A(ram[2524]), .B(n12878), .Y(n2751) );
  OAI21X1 U5256 ( .A(n12696), .B(n12878), .C(n2752), .Y(n6962) );
  NAND2X1 U5257 ( .A(ram[2525]), .B(n12878), .Y(n2752) );
  OAI21X1 U5258 ( .A(n12691), .B(n12878), .C(n2753), .Y(n6963) );
  NAND2X1 U5259 ( .A(ram[2526]), .B(n12878), .Y(n2753) );
  OAI21X1 U5260 ( .A(n12685), .B(n12878), .C(n2754), .Y(n6964) );
  NAND2X1 U5261 ( .A(ram[2527]), .B(n12878), .Y(n2754) );
  OAI21X1 U5263 ( .A(n12775), .B(n12877), .C(n2756), .Y(n6965) );
  NAND2X1 U5264 ( .A(ram[2528]), .B(n12877), .Y(n2756) );
  OAI21X1 U5265 ( .A(n12769), .B(n12877), .C(n2757), .Y(n6966) );
  NAND2X1 U5266 ( .A(ram[2529]), .B(n12877), .Y(n2757) );
  OAI21X1 U5267 ( .A(n12762), .B(n12877), .C(n2758), .Y(n6967) );
  NAND2X1 U5268 ( .A(ram[2530]), .B(n12877), .Y(n2758) );
  OAI21X1 U5269 ( .A(n12756), .B(n12877), .C(n2759), .Y(n6968) );
  NAND2X1 U5270 ( .A(ram[2531]), .B(n12877), .Y(n2759) );
  OAI21X1 U5271 ( .A(n12750), .B(n12877), .C(n2760), .Y(n6969) );
  NAND2X1 U5272 ( .A(ram[2532]), .B(n12877), .Y(n2760) );
  OAI21X1 U5273 ( .A(n12744), .B(n12877), .C(n2761), .Y(n6970) );
  NAND2X1 U5274 ( .A(ram[2533]), .B(n12877), .Y(n2761) );
  OAI21X1 U5275 ( .A(n12738), .B(n12877), .C(n2762), .Y(n6971) );
  NAND2X1 U5276 ( .A(ram[2534]), .B(n12877), .Y(n2762) );
  OAI21X1 U5277 ( .A(n12732), .B(n12877), .C(n2763), .Y(n6972) );
  NAND2X1 U5278 ( .A(ram[2535]), .B(n12877), .Y(n2763) );
  OAI21X1 U5279 ( .A(n12726), .B(n12877), .C(n2764), .Y(n6973) );
  NAND2X1 U5280 ( .A(ram[2536]), .B(n12877), .Y(n2764) );
  OAI21X1 U5281 ( .A(n12720), .B(n12877), .C(n2765), .Y(n6974) );
  NAND2X1 U5282 ( .A(ram[2537]), .B(n12877), .Y(n2765) );
  OAI21X1 U5283 ( .A(n12714), .B(n12877), .C(n2766), .Y(n6975) );
  NAND2X1 U5284 ( .A(ram[2538]), .B(n12877), .Y(n2766) );
  OAI21X1 U5285 ( .A(n12708), .B(n12877), .C(n2767), .Y(n6976) );
  NAND2X1 U5286 ( .A(ram[2539]), .B(n12877), .Y(n2767) );
  OAI21X1 U5287 ( .A(n12702), .B(n12877), .C(n2768), .Y(n6977) );
  NAND2X1 U5288 ( .A(ram[2540]), .B(n12877), .Y(n2768) );
  OAI21X1 U5289 ( .A(n12696), .B(n12877), .C(n2769), .Y(n6978) );
  NAND2X1 U5290 ( .A(ram[2541]), .B(n12877), .Y(n2769) );
  OAI21X1 U5291 ( .A(n12691), .B(n12877), .C(n2770), .Y(n6979) );
  NAND2X1 U5292 ( .A(ram[2542]), .B(n12877), .Y(n2770) );
  OAI21X1 U5293 ( .A(n12685), .B(n12877), .C(n2771), .Y(n6980) );
  NAND2X1 U5294 ( .A(ram[2543]), .B(n12877), .Y(n2771) );
  OAI21X1 U5296 ( .A(n12774), .B(n12876), .C(n2773), .Y(n6981) );
  NAND2X1 U5297 ( .A(ram[2544]), .B(n12876), .Y(n2773) );
  OAI21X1 U5298 ( .A(n12768), .B(n12876), .C(n2774), .Y(n6982) );
  NAND2X1 U5299 ( .A(ram[2545]), .B(n12876), .Y(n2774) );
  OAI21X1 U5300 ( .A(n12763), .B(n12876), .C(n2775), .Y(n6983) );
  NAND2X1 U5301 ( .A(ram[2546]), .B(n12876), .Y(n2775) );
  OAI21X1 U5302 ( .A(n12757), .B(n12876), .C(n2776), .Y(n6984) );
  NAND2X1 U5303 ( .A(ram[2547]), .B(n12876), .Y(n2776) );
  OAI21X1 U5304 ( .A(n12751), .B(n12876), .C(n2777), .Y(n6985) );
  NAND2X1 U5305 ( .A(ram[2548]), .B(n12876), .Y(n2777) );
  OAI21X1 U5306 ( .A(n12745), .B(n12876), .C(n2778), .Y(n6986) );
  NAND2X1 U5307 ( .A(ram[2549]), .B(n12876), .Y(n2778) );
  OAI21X1 U5308 ( .A(n12739), .B(n12876), .C(n2779), .Y(n6987) );
  NAND2X1 U5309 ( .A(ram[2550]), .B(n12876), .Y(n2779) );
  OAI21X1 U5310 ( .A(n12733), .B(n12876), .C(n2780), .Y(n6988) );
  NAND2X1 U5311 ( .A(ram[2551]), .B(n12876), .Y(n2780) );
  OAI21X1 U5312 ( .A(n12727), .B(n12876), .C(n2781), .Y(n6989) );
  NAND2X1 U5313 ( .A(ram[2552]), .B(n12876), .Y(n2781) );
  OAI21X1 U5314 ( .A(n12721), .B(n12876), .C(n2782), .Y(n6990) );
  NAND2X1 U5315 ( .A(ram[2553]), .B(n12876), .Y(n2782) );
  OAI21X1 U5316 ( .A(n12715), .B(n12876), .C(n2783), .Y(n6991) );
  NAND2X1 U5317 ( .A(ram[2554]), .B(n12876), .Y(n2783) );
  OAI21X1 U5318 ( .A(n12709), .B(n12876), .C(n2784), .Y(n6992) );
  NAND2X1 U5319 ( .A(ram[2555]), .B(n12876), .Y(n2784) );
  OAI21X1 U5320 ( .A(n12703), .B(n12876), .C(n2785), .Y(n6993) );
  NAND2X1 U5321 ( .A(ram[2556]), .B(n12876), .Y(n2785) );
  OAI21X1 U5322 ( .A(n12697), .B(n12876), .C(n2786), .Y(n6994) );
  NAND2X1 U5323 ( .A(ram[2557]), .B(n12876), .Y(n2786) );
  OAI21X1 U5324 ( .A(n12690), .B(n12876), .C(n2787), .Y(n6995) );
  NAND2X1 U5325 ( .A(ram[2558]), .B(n12876), .Y(n2787) );
  OAI21X1 U5326 ( .A(n12684), .B(n12876), .C(n2788), .Y(n6996) );
  NAND2X1 U5327 ( .A(ram[2559]), .B(n12876), .Y(n2788) );
  NAND3X1 U5329 ( .A(n601), .B(mem_write_en), .C(n2516), .Y(n2789) );
  OAI21X1 U5330 ( .A(n12775), .B(n12875), .C(n2791), .Y(n6997) );
  NAND2X1 U5331 ( .A(ram[2560]), .B(n12875), .Y(n2791) );
  OAI21X1 U5332 ( .A(n12769), .B(n12875), .C(n2792), .Y(n6998) );
  NAND2X1 U5333 ( .A(ram[2561]), .B(n12875), .Y(n2792) );
  OAI21X1 U5334 ( .A(n12765), .B(n12875), .C(n2793), .Y(n6999) );
  NAND2X1 U5335 ( .A(ram[2562]), .B(n12875), .Y(n2793) );
  OAI21X1 U5336 ( .A(n12759), .B(n12875), .C(n2794), .Y(n7000) );
  NAND2X1 U5337 ( .A(ram[2563]), .B(n12875), .Y(n2794) );
  OAI21X1 U5338 ( .A(n12753), .B(n12875), .C(n2795), .Y(n7001) );
  NAND2X1 U5339 ( .A(ram[2564]), .B(n12875), .Y(n2795) );
  OAI21X1 U5340 ( .A(n12747), .B(n12875), .C(n2796), .Y(n7002) );
  NAND2X1 U5341 ( .A(ram[2565]), .B(n12875), .Y(n2796) );
  OAI21X1 U5342 ( .A(n12741), .B(n12875), .C(n2797), .Y(n7003) );
  NAND2X1 U5343 ( .A(ram[2566]), .B(n12875), .Y(n2797) );
  OAI21X1 U5344 ( .A(n12735), .B(n12875), .C(n2798), .Y(n7004) );
  NAND2X1 U5345 ( .A(ram[2567]), .B(n12875), .Y(n2798) );
  OAI21X1 U5346 ( .A(n12729), .B(n12875), .C(n2799), .Y(n7005) );
  NAND2X1 U5347 ( .A(ram[2568]), .B(n12875), .Y(n2799) );
  OAI21X1 U5348 ( .A(n12723), .B(n12875), .C(n2800), .Y(n7006) );
  NAND2X1 U5349 ( .A(ram[2569]), .B(n12875), .Y(n2800) );
  OAI21X1 U5350 ( .A(n12717), .B(n12875), .C(n2801), .Y(n7007) );
  NAND2X1 U5351 ( .A(ram[2570]), .B(n12875), .Y(n2801) );
  OAI21X1 U5352 ( .A(n12711), .B(n12875), .C(n2802), .Y(n7008) );
  NAND2X1 U5353 ( .A(ram[2571]), .B(n12875), .Y(n2802) );
  OAI21X1 U5354 ( .A(n12705), .B(n12875), .C(n2803), .Y(n7009) );
  NAND2X1 U5355 ( .A(ram[2572]), .B(n12875), .Y(n2803) );
  OAI21X1 U5356 ( .A(n12699), .B(n12875), .C(n2804), .Y(n7010) );
  NAND2X1 U5357 ( .A(ram[2573]), .B(n12875), .Y(n2804) );
  OAI21X1 U5358 ( .A(n12691), .B(n12875), .C(n2805), .Y(n7011) );
  NAND2X1 U5359 ( .A(ram[2574]), .B(n12875), .Y(n2805) );
  OAI21X1 U5360 ( .A(n12685), .B(n12875), .C(n2806), .Y(n7012) );
  NAND2X1 U5361 ( .A(ram[2575]), .B(n12875), .Y(n2806) );
  OAI21X1 U5363 ( .A(n12774), .B(n12874), .C(n2808), .Y(n7013) );
  NAND2X1 U5364 ( .A(ram[2576]), .B(n12874), .Y(n2808) );
  OAI21X1 U5365 ( .A(n12768), .B(n12874), .C(n2809), .Y(n7014) );
  NAND2X1 U5366 ( .A(ram[2577]), .B(n12874), .Y(n2809) );
  OAI21X1 U5367 ( .A(n12765), .B(n12874), .C(n2810), .Y(n7015) );
  NAND2X1 U5368 ( .A(ram[2578]), .B(n12874), .Y(n2810) );
  OAI21X1 U5369 ( .A(n12759), .B(n12874), .C(n2811), .Y(n7016) );
  NAND2X1 U5370 ( .A(ram[2579]), .B(n12874), .Y(n2811) );
  OAI21X1 U5371 ( .A(n12753), .B(n12874), .C(n2812), .Y(n7017) );
  NAND2X1 U5372 ( .A(ram[2580]), .B(n12874), .Y(n2812) );
  OAI21X1 U5373 ( .A(n12747), .B(n12874), .C(n2813), .Y(n7018) );
  NAND2X1 U5374 ( .A(ram[2581]), .B(n12874), .Y(n2813) );
  OAI21X1 U5375 ( .A(n12741), .B(n12874), .C(n2814), .Y(n7019) );
  NAND2X1 U5376 ( .A(ram[2582]), .B(n12874), .Y(n2814) );
  OAI21X1 U5377 ( .A(n12735), .B(n12874), .C(n2815), .Y(n7020) );
  NAND2X1 U5378 ( .A(ram[2583]), .B(n12874), .Y(n2815) );
  OAI21X1 U5379 ( .A(n12729), .B(n12874), .C(n2816), .Y(n7021) );
  NAND2X1 U5380 ( .A(ram[2584]), .B(n12874), .Y(n2816) );
  OAI21X1 U5381 ( .A(n12723), .B(n12874), .C(n2817), .Y(n7022) );
  NAND2X1 U5382 ( .A(ram[2585]), .B(n12874), .Y(n2817) );
  OAI21X1 U5383 ( .A(n12717), .B(n12874), .C(n2818), .Y(n7023) );
  NAND2X1 U5384 ( .A(ram[2586]), .B(n12874), .Y(n2818) );
  OAI21X1 U5385 ( .A(n12711), .B(n12874), .C(n2819), .Y(n7024) );
  NAND2X1 U5386 ( .A(ram[2587]), .B(n12874), .Y(n2819) );
  OAI21X1 U5387 ( .A(n12705), .B(n12874), .C(n2820), .Y(n7025) );
  NAND2X1 U5388 ( .A(ram[2588]), .B(n12874), .Y(n2820) );
  OAI21X1 U5389 ( .A(n12699), .B(n12874), .C(n2821), .Y(n7026) );
  NAND2X1 U5390 ( .A(ram[2589]), .B(n12874), .Y(n2821) );
  OAI21X1 U5391 ( .A(n12690), .B(n12874), .C(n2822), .Y(n7027) );
  NAND2X1 U5392 ( .A(ram[2590]), .B(n12874), .Y(n2822) );
  OAI21X1 U5393 ( .A(n12684), .B(n12874), .C(n2823), .Y(n7028) );
  NAND2X1 U5394 ( .A(ram[2591]), .B(n12874), .Y(n2823) );
  OAI21X1 U5396 ( .A(n12776), .B(n12873), .C(n2825), .Y(n7029) );
  NAND2X1 U5397 ( .A(ram[2592]), .B(n12873), .Y(n2825) );
  OAI21X1 U5398 ( .A(n12770), .B(n12873), .C(n2826), .Y(n7030) );
  NAND2X1 U5399 ( .A(ram[2593]), .B(n12873), .Y(n2826) );
  OAI21X1 U5400 ( .A(n12765), .B(n12873), .C(n2827), .Y(n7031) );
  NAND2X1 U5401 ( .A(ram[2594]), .B(n12873), .Y(n2827) );
  OAI21X1 U5402 ( .A(n12759), .B(n12873), .C(n2828), .Y(n7032) );
  NAND2X1 U5403 ( .A(ram[2595]), .B(n12873), .Y(n2828) );
  OAI21X1 U5404 ( .A(n12753), .B(n12873), .C(n2829), .Y(n7033) );
  NAND2X1 U5405 ( .A(ram[2596]), .B(n12873), .Y(n2829) );
  OAI21X1 U5406 ( .A(n12747), .B(n12873), .C(n2830), .Y(n7034) );
  NAND2X1 U5407 ( .A(ram[2597]), .B(n12873), .Y(n2830) );
  OAI21X1 U5408 ( .A(n12741), .B(n12873), .C(n2831), .Y(n7035) );
  NAND2X1 U5409 ( .A(ram[2598]), .B(n12873), .Y(n2831) );
  OAI21X1 U5410 ( .A(n12735), .B(n12873), .C(n2832), .Y(n7036) );
  NAND2X1 U5411 ( .A(ram[2599]), .B(n12873), .Y(n2832) );
  OAI21X1 U5412 ( .A(n12729), .B(n12873), .C(n2833), .Y(n7037) );
  NAND2X1 U5413 ( .A(ram[2600]), .B(n12873), .Y(n2833) );
  OAI21X1 U5414 ( .A(n12723), .B(n12873), .C(n2834), .Y(n7038) );
  NAND2X1 U5415 ( .A(ram[2601]), .B(n12873), .Y(n2834) );
  OAI21X1 U5416 ( .A(n12717), .B(n12873), .C(n2835), .Y(n7039) );
  NAND2X1 U5417 ( .A(ram[2602]), .B(n12873), .Y(n2835) );
  OAI21X1 U5418 ( .A(n12711), .B(n12873), .C(n2836), .Y(n7040) );
  NAND2X1 U5419 ( .A(ram[2603]), .B(n12873), .Y(n2836) );
  OAI21X1 U5420 ( .A(n12705), .B(n12873), .C(n2837), .Y(n7041) );
  NAND2X1 U5421 ( .A(ram[2604]), .B(n12873), .Y(n2837) );
  OAI21X1 U5422 ( .A(n12699), .B(n12873), .C(n2838), .Y(n7042) );
  NAND2X1 U5423 ( .A(ram[2605]), .B(n12873), .Y(n2838) );
  OAI21X1 U5424 ( .A(n12692), .B(n12873), .C(n2839), .Y(n7043) );
  NAND2X1 U5425 ( .A(ram[2606]), .B(n12873), .Y(n2839) );
  OAI21X1 U5426 ( .A(n12686), .B(n12873), .C(n2840), .Y(n7044) );
  NAND2X1 U5427 ( .A(ram[2607]), .B(n12873), .Y(n2840) );
  OAI21X1 U5429 ( .A(n12779), .B(n12872), .C(n2842), .Y(n7045) );
  NAND2X1 U5430 ( .A(ram[2608]), .B(n12872), .Y(n2842) );
  OAI21X1 U5431 ( .A(n12773), .B(n12872), .C(n2843), .Y(n7046) );
  NAND2X1 U5432 ( .A(ram[2609]), .B(n12872), .Y(n2843) );
  OAI21X1 U5433 ( .A(n12767), .B(n12872), .C(n2844), .Y(n7047) );
  NAND2X1 U5434 ( .A(ram[2610]), .B(n12872), .Y(n2844) );
  OAI21X1 U5435 ( .A(n12761), .B(n12872), .C(n2845), .Y(n7048) );
  NAND2X1 U5436 ( .A(ram[2611]), .B(n12872), .Y(n2845) );
  OAI21X1 U5437 ( .A(n12755), .B(n12872), .C(n2846), .Y(n7049) );
  NAND2X1 U5438 ( .A(ram[2612]), .B(n12872), .Y(n2846) );
  OAI21X1 U5439 ( .A(n12749), .B(n12872), .C(n2847), .Y(n7050) );
  NAND2X1 U5440 ( .A(ram[2613]), .B(n12872), .Y(n2847) );
  OAI21X1 U5441 ( .A(n12743), .B(n12872), .C(n2848), .Y(n7051) );
  NAND2X1 U5442 ( .A(ram[2614]), .B(n12872), .Y(n2848) );
  OAI21X1 U5443 ( .A(n12737), .B(n12872), .C(n2849), .Y(n7052) );
  NAND2X1 U5444 ( .A(ram[2615]), .B(n12872), .Y(n2849) );
  OAI21X1 U5445 ( .A(n12731), .B(n12872), .C(n2850), .Y(n7053) );
  NAND2X1 U5446 ( .A(ram[2616]), .B(n12872), .Y(n2850) );
  OAI21X1 U5447 ( .A(n12725), .B(n12872), .C(n2851), .Y(n7054) );
  NAND2X1 U5448 ( .A(ram[2617]), .B(n12872), .Y(n2851) );
  OAI21X1 U5449 ( .A(n12719), .B(n12872), .C(n2852), .Y(n7055) );
  NAND2X1 U5450 ( .A(ram[2618]), .B(n12872), .Y(n2852) );
  OAI21X1 U5451 ( .A(n12713), .B(n12872), .C(n2853), .Y(n7056) );
  NAND2X1 U5452 ( .A(ram[2619]), .B(n12872), .Y(n2853) );
  OAI21X1 U5453 ( .A(n12707), .B(n12872), .C(n2854), .Y(n7057) );
  NAND2X1 U5454 ( .A(ram[2620]), .B(n12872), .Y(n2854) );
  OAI21X1 U5455 ( .A(n12701), .B(n12872), .C(n2855), .Y(n7058) );
  NAND2X1 U5456 ( .A(ram[2621]), .B(n12872), .Y(n2855) );
  OAI21X1 U5457 ( .A(n12695), .B(n12872), .C(n2856), .Y(n7059) );
  NAND2X1 U5458 ( .A(ram[2622]), .B(n12872), .Y(n2856) );
  OAI21X1 U5459 ( .A(n12689), .B(n12872), .C(n2857), .Y(n7060) );
  NAND2X1 U5460 ( .A(ram[2623]), .B(n12872), .Y(n2857) );
  OAI21X1 U5462 ( .A(n12778), .B(n12871), .C(n2859), .Y(n7061) );
  NAND2X1 U5463 ( .A(ram[2624]), .B(n12871), .Y(n2859) );
  OAI21X1 U5464 ( .A(n12772), .B(n12871), .C(n2860), .Y(n7062) );
  NAND2X1 U5465 ( .A(ram[2625]), .B(n12871), .Y(n2860) );
  OAI21X1 U5466 ( .A(n12766), .B(n12871), .C(n2861), .Y(n7063) );
  NAND2X1 U5467 ( .A(ram[2626]), .B(n12871), .Y(n2861) );
  OAI21X1 U5468 ( .A(n12760), .B(n12871), .C(n2862), .Y(n7064) );
  NAND2X1 U5469 ( .A(ram[2627]), .B(n12871), .Y(n2862) );
  OAI21X1 U5470 ( .A(n12754), .B(n12871), .C(n2863), .Y(n7065) );
  NAND2X1 U5471 ( .A(ram[2628]), .B(n12871), .Y(n2863) );
  OAI21X1 U5472 ( .A(n12748), .B(n12871), .C(n2864), .Y(n7066) );
  NAND2X1 U5473 ( .A(ram[2629]), .B(n12871), .Y(n2864) );
  OAI21X1 U5474 ( .A(n12742), .B(n12871), .C(n2865), .Y(n7067) );
  NAND2X1 U5475 ( .A(ram[2630]), .B(n12871), .Y(n2865) );
  OAI21X1 U5476 ( .A(n12736), .B(n12871), .C(n2866), .Y(n7068) );
  NAND2X1 U5477 ( .A(ram[2631]), .B(n12871), .Y(n2866) );
  OAI21X1 U5478 ( .A(n12730), .B(n12871), .C(n2867), .Y(n7069) );
  NAND2X1 U5479 ( .A(ram[2632]), .B(n12871), .Y(n2867) );
  OAI21X1 U5480 ( .A(n12724), .B(n12871), .C(n2868), .Y(n7070) );
  NAND2X1 U5481 ( .A(ram[2633]), .B(n12871), .Y(n2868) );
  OAI21X1 U5482 ( .A(n12718), .B(n12871), .C(n2869), .Y(n7071) );
  NAND2X1 U5483 ( .A(ram[2634]), .B(n12871), .Y(n2869) );
  OAI21X1 U5484 ( .A(n12712), .B(n12871), .C(n2870), .Y(n7072) );
  NAND2X1 U5485 ( .A(ram[2635]), .B(n12871), .Y(n2870) );
  OAI21X1 U5486 ( .A(n12706), .B(n12871), .C(n2871), .Y(n7073) );
  NAND2X1 U5487 ( .A(ram[2636]), .B(n12871), .Y(n2871) );
  OAI21X1 U5488 ( .A(n12700), .B(n12871), .C(n2872), .Y(n7074) );
  NAND2X1 U5489 ( .A(ram[2637]), .B(n12871), .Y(n2872) );
  OAI21X1 U5490 ( .A(n12694), .B(n12871), .C(n2873), .Y(n7075) );
  NAND2X1 U5491 ( .A(ram[2638]), .B(n12871), .Y(n2873) );
  OAI21X1 U5492 ( .A(n12688), .B(n12871), .C(n2874), .Y(n7076) );
  NAND2X1 U5493 ( .A(ram[2639]), .B(n12871), .Y(n2874) );
  OAI21X1 U5495 ( .A(n12777), .B(n12870), .C(n2876), .Y(n7077) );
  NAND2X1 U5496 ( .A(ram[2640]), .B(n12870), .Y(n2876) );
  OAI21X1 U5497 ( .A(n12771), .B(n12870), .C(n2877), .Y(n7078) );
  NAND2X1 U5498 ( .A(ram[2641]), .B(n12870), .Y(n2877) );
  OAI21X1 U5499 ( .A(n12765), .B(n12870), .C(n2878), .Y(n7079) );
  NAND2X1 U5500 ( .A(ram[2642]), .B(n12870), .Y(n2878) );
  OAI21X1 U5501 ( .A(n12759), .B(n12870), .C(n2879), .Y(n7080) );
  NAND2X1 U5502 ( .A(ram[2643]), .B(n12870), .Y(n2879) );
  OAI21X1 U5503 ( .A(n12753), .B(n12870), .C(n2880), .Y(n7081) );
  NAND2X1 U5504 ( .A(ram[2644]), .B(n12870), .Y(n2880) );
  OAI21X1 U5505 ( .A(n12747), .B(n12870), .C(n2881), .Y(n7082) );
  NAND2X1 U5506 ( .A(ram[2645]), .B(n12870), .Y(n2881) );
  OAI21X1 U5507 ( .A(n12741), .B(n12870), .C(n2882), .Y(n7083) );
  NAND2X1 U5508 ( .A(ram[2646]), .B(n12870), .Y(n2882) );
  OAI21X1 U5509 ( .A(n12735), .B(n12870), .C(n2883), .Y(n7084) );
  NAND2X1 U5510 ( .A(ram[2647]), .B(n12870), .Y(n2883) );
  OAI21X1 U5511 ( .A(n12729), .B(n12870), .C(n2884), .Y(n7085) );
  NAND2X1 U5512 ( .A(ram[2648]), .B(n12870), .Y(n2884) );
  OAI21X1 U5513 ( .A(n12723), .B(n12870), .C(n2885), .Y(n7086) );
  NAND2X1 U5514 ( .A(ram[2649]), .B(n12870), .Y(n2885) );
  OAI21X1 U5515 ( .A(n12717), .B(n12870), .C(n2886), .Y(n7087) );
  NAND2X1 U5516 ( .A(ram[2650]), .B(n12870), .Y(n2886) );
  OAI21X1 U5517 ( .A(n12711), .B(n12870), .C(n2887), .Y(n7088) );
  NAND2X1 U5518 ( .A(ram[2651]), .B(n12870), .Y(n2887) );
  OAI21X1 U5519 ( .A(n12705), .B(n12870), .C(n2888), .Y(n7089) );
  NAND2X1 U5520 ( .A(ram[2652]), .B(n12870), .Y(n2888) );
  OAI21X1 U5521 ( .A(n12699), .B(n12870), .C(n2889), .Y(n7090) );
  NAND2X1 U5522 ( .A(ram[2653]), .B(n12870), .Y(n2889) );
  OAI21X1 U5523 ( .A(n12693), .B(n12870), .C(n2890), .Y(n7091) );
  NAND2X1 U5524 ( .A(ram[2654]), .B(n12870), .Y(n2890) );
  OAI21X1 U5525 ( .A(n12687), .B(n12870), .C(n2891), .Y(n7092) );
  NAND2X1 U5526 ( .A(ram[2655]), .B(n12870), .Y(n2891) );
  OAI21X1 U5528 ( .A(n12776), .B(n12869), .C(n2893), .Y(n7093) );
  NAND2X1 U5529 ( .A(ram[2656]), .B(n12869), .Y(n2893) );
  OAI21X1 U5530 ( .A(n12770), .B(n12869), .C(n2894), .Y(n7094) );
  NAND2X1 U5531 ( .A(ram[2657]), .B(n12869), .Y(n2894) );
  OAI21X1 U5532 ( .A(n12763), .B(n12869), .C(n2895), .Y(n7095) );
  NAND2X1 U5533 ( .A(ram[2658]), .B(n12869), .Y(n2895) );
  OAI21X1 U5534 ( .A(n12757), .B(n12869), .C(n2896), .Y(n7096) );
  NAND2X1 U5535 ( .A(ram[2659]), .B(n12869), .Y(n2896) );
  OAI21X1 U5536 ( .A(n12751), .B(n12869), .C(n2897), .Y(n7097) );
  NAND2X1 U5537 ( .A(ram[2660]), .B(n12869), .Y(n2897) );
  OAI21X1 U5538 ( .A(n12745), .B(n12869), .C(n2898), .Y(n7098) );
  NAND2X1 U5539 ( .A(ram[2661]), .B(n12869), .Y(n2898) );
  OAI21X1 U5540 ( .A(n12739), .B(n12869), .C(n2899), .Y(n7099) );
  NAND2X1 U5541 ( .A(ram[2662]), .B(n12869), .Y(n2899) );
  OAI21X1 U5542 ( .A(n12733), .B(n12869), .C(n2900), .Y(n7100) );
  NAND2X1 U5543 ( .A(ram[2663]), .B(n12869), .Y(n2900) );
  OAI21X1 U5544 ( .A(n12727), .B(n12869), .C(n2901), .Y(n7101) );
  NAND2X1 U5545 ( .A(ram[2664]), .B(n12869), .Y(n2901) );
  OAI21X1 U5546 ( .A(n12721), .B(n12869), .C(n2902), .Y(n7102) );
  NAND2X1 U5547 ( .A(ram[2665]), .B(n12869), .Y(n2902) );
  OAI21X1 U5548 ( .A(n12715), .B(n12869), .C(n2903), .Y(n7103) );
  NAND2X1 U5549 ( .A(ram[2666]), .B(n12869), .Y(n2903) );
  OAI21X1 U5550 ( .A(n12709), .B(n12869), .C(n2904), .Y(n7104) );
  NAND2X1 U5551 ( .A(ram[2667]), .B(n12869), .Y(n2904) );
  OAI21X1 U5552 ( .A(n12703), .B(n12869), .C(n2905), .Y(n7105) );
  NAND2X1 U5553 ( .A(ram[2668]), .B(n12869), .Y(n2905) );
  OAI21X1 U5554 ( .A(n12697), .B(n12869), .C(n2906), .Y(n7106) );
  NAND2X1 U5555 ( .A(ram[2669]), .B(n12869), .Y(n2906) );
  OAI21X1 U5556 ( .A(n12692), .B(n12869), .C(n2907), .Y(n7107) );
  NAND2X1 U5557 ( .A(ram[2670]), .B(n12869), .Y(n2907) );
  OAI21X1 U5558 ( .A(n12686), .B(n12869), .C(n2908), .Y(n7108) );
  NAND2X1 U5559 ( .A(ram[2671]), .B(n12869), .Y(n2908) );
  OAI21X1 U5561 ( .A(n12776), .B(n12868), .C(n2910), .Y(n7109) );
  NAND2X1 U5562 ( .A(ram[2672]), .B(n12868), .Y(n2910) );
  OAI21X1 U5563 ( .A(n12770), .B(n12868), .C(n2911), .Y(n7110) );
  NAND2X1 U5564 ( .A(ram[2673]), .B(n12868), .Y(n2911) );
  OAI21X1 U5565 ( .A(n12764), .B(n12868), .C(n2912), .Y(n7111) );
  NAND2X1 U5566 ( .A(ram[2674]), .B(n12868), .Y(n2912) );
  OAI21X1 U5567 ( .A(n12758), .B(n12868), .C(n2913), .Y(n7112) );
  NAND2X1 U5568 ( .A(ram[2675]), .B(n12868), .Y(n2913) );
  OAI21X1 U5569 ( .A(n12752), .B(n12868), .C(n2914), .Y(n7113) );
  NAND2X1 U5570 ( .A(ram[2676]), .B(n12868), .Y(n2914) );
  OAI21X1 U5571 ( .A(n12746), .B(n12868), .C(n2915), .Y(n7114) );
  NAND2X1 U5572 ( .A(ram[2677]), .B(n12868), .Y(n2915) );
  OAI21X1 U5573 ( .A(n12740), .B(n12868), .C(n2916), .Y(n7115) );
  NAND2X1 U5574 ( .A(ram[2678]), .B(n12868), .Y(n2916) );
  OAI21X1 U5575 ( .A(n12734), .B(n12868), .C(n2917), .Y(n7116) );
  NAND2X1 U5576 ( .A(ram[2679]), .B(n12868), .Y(n2917) );
  OAI21X1 U5577 ( .A(n12728), .B(n12868), .C(n2918), .Y(n7117) );
  NAND2X1 U5578 ( .A(ram[2680]), .B(n12868), .Y(n2918) );
  OAI21X1 U5579 ( .A(n12722), .B(n12868), .C(n2919), .Y(n7118) );
  NAND2X1 U5580 ( .A(ram[2681]), .B(n12868), .Y(n2919) );
  OAI21X1 U5581 ( .A(n12716), .B(n12868), .C(n2920), .Y(n7119) );
  NAND2X1 U5582 ( .A(ram[2682]), .B(n12868), .Y(n2920) );
  OAI21X1 U5583 ( .A(n12710), .B(n12868), .C(n2921), .Y(n7120) );
  NAND2X1 U5584 ( .A(ram[2683]), .B(n12868), .Y(n2921) );
  OAI21X1 U5585 ( .A(n12704), .B(n12868), .C(n2922), .Y(n7121) );
  NAND2X1 U5586 ( .A(ram[2684]), .B(n12868), .Y(n2922) );
  OAI21X1 U5587 ( .A(n12698), .B(n12868), .C(n2923), .Y(n7122) );
  NAND2X1 U5588 ( .A(ram[2685]), .B(n12868), .Y(n2923) );
  OAI21X1 U5589 ( .A(n12692), .B(n12868), .C(n2924), .Y(n7123) );
  NAND2X1 U5590 ( .A(ram[2686]), .B(n12868), .Y(n2924) );
  OAI21X1 U5591 ( .A(n12686), .B(n12868), .C(n2925), .Y(n7124) );
  NAND2X1 U5592 ( .A(ram[2687]), .B(n12868), .Y(n2925) );
  OAI21X1 U5594 ( .A(n12776), .B(n12867), .C(n2927), .Y(n7125) );
  NAND2X1 U5595 ( .A(ram[2688]), .B(n12867), .Y(n2927) );
  OAI21X1 U5596 ( .A(n12770), .B(n12867), .C(n2928), .Y(n7126) );
  NAND2X1 U5597 ( .A(ram[2689]), .B(n12867), .Y(n2928) );
  OAI21X1 U5598 ( .A(n12764), .B(n12867), .C(n2929), .Y(n7127) );
  NAND2X1 U5599 ( .A(ram[2690]), .B(n12867), .Y(n2929) );
  OAI21X1 U5600 ( .A(n12758), .B(n12867), .C(n2930), .Y(n7128) );
  NAND2X1 U5601 ( .A(ram[2691]), .B(n12867), .Y(n2930) );
  OAI21X1 U5602 ( .A(n12752), .B(n12867), .C(n2931), .Y(n7129) );
  NAND2X1 U5603 ( .A(ram[2692]), .B(n12867), .Y(n2931) );
  OAI21X1 U5604 ( .A(n12746), .B(n12867), .C(n2932), .Y(n7130) );
  NAND2X1 U5605 ( .A(ram[2693]), .B(n12867), .Y(n2932) );
  OAI21X1 U5606 ( .A(n12740), .B(n12867), .C(n2933), .Y(n7131) );
  NAND2X1 U5607 ( .A(ram[2694]), .B(n12867), .Y(n2933) );
  OAI21X1 U5608 ( .A(n12734), .B(n12867), .C(n2934), .Y(n7132) );
  NAND2X1 U5609 ( .A(ram[2695]), .B(n12867), .Y(n2934) );
  OAI21X1 U5610 ( .A(n12728), .B(n12867), .C(n2935), .Y(n7133) );
  NAND2X1 U5611 ( .A(ram[2696]), .B(n12867), .Y(n2935) );
  OAI21X1 U5612 ( .A(n12722), .B(n12867), .C(n2936), .Y(n7134) );
  NAND2X1 U5613 ( .A(ram[2697]), .B(n12867), .Y(n2936) );
  OAI21X1 U5614 ( .A(n12716), .B(n12867), .C(n2937), .Y(n7135) );
  NAND2X1 U5615 ( .A(ram[2698]), .B(n12867), .Y(n2937) );
  OAI21X1 U5616 ( .A(n12710), .B(n12867), .C(n2938), .Y(n7136) );
  NAND2X1 U5617 ( .A(ram[2699]), .B(n12867), .Y(n2938) );
  OAI21X1 U5618 ( .A(n12704), .B(n12867), .C(n2939), .Y(n7137) );
  NAND2X1 U5619 ( .A(ram[2700]), .B(n12867), .Y(n2939) );
  OAI21X1 U5620 ( .A(n12698), .B(n12867), .C(n2940), .Y(n7138) );
  NAND2X1 U5621 ( .A(ram[2701]), .B(n12867), .Y(n2940) );
  OAI21X1 U5622 ( .A(n12692), .B(n12867), .C(n2941), .Y(n7139) );
  NAND2X1 U5623 ( .A(ram[2702]), .B(n12867), .Y(n2941) );
  OAI21X1 U5624 ( .A(n12686), .B(n12867), .C(n2942), .Y(n7140) );
  NAND2X1 U5625 ( .A(ram[2703]), .B(n12867), .Y(n2942) );
  OAI21X1 U5627 ( .A(n12779), .B(n12866), .C(n2944), .Y(n7141) );
  NAND2X1 U5628 ( .A(ram[2704]), .B(n12866), .Y(n2944) );
  OAI21X1 U5629 ( .A(n12773), .B(n12866), .C(n2945), .Y(n7142) );
  NAND2X1 U5630 ( .A(ram[2705]), .B(n12866), .Y(n2945) );
  OAI21X1 U5631 ( .A(n12764), .B(n12866), .C(n2946), .Y(n7143) );
  NAND2X1 U5632 ( .A(ram[2706]), .B(n12866), .Y(n2946) );
  OAI21X1 U5633 ( .A(n12758), .B(n12866), .C(n2947), .Y(n7144) );
  NAND2X1 U5634 ( .A(ram[2707]), .B(n12866), .Y(n2947) );
  OAI21X1 U5635 ( .A(n12752), .B(n12866), .C(n2948), .Y(n7145) );
  NAND2X1 U5636 ( .A(ram[2708]), .B(n12866), .Y(n2948) );
  OAI21X1 U5637 ( .A(n12746), .B(n12866), .C(n2949), .Y(n7146) );
  NAND2X1 U5638 ( .A(ram[2709]), .B(n12866), .Y(n2949) );
  OAI21X1 U5639 ( .A(n12740), .B(n12866), .C(n2950), .Y(n7147) );
  NAND2X1 U5640 ( .A(ram[2710]), .B(n12866), .Y(n2950) );
  OAI21X1 U5641 ( .A(n12734), .B(n12866), .C(n2951), .Y(n7148) );
  NAND2X1 U5642 ( .A(ram[2711]), .B(n12866), .Y(n2951) );
  OAI21X1 U5643 ( .A(n12728), .B(n12866), .C(n2952), .Y(n7149) );
  NAND2X1 U5644 ( .A(ram[2712]), .B(n12866), .Y(n2952) );
  OAI21X1 U5645 ( .A(n12722), .B(n12866), .C(n2953), .Y(n7150) );
  NAND2X1 U5646 ( .A(ram[2713]), .B(n12866), .Y(n2953) );
  OAI21X1 U5647 ( .A(n12716), .B(n12866), .C(n2954), .Y(n7151) );
  NAND2X1 U5648 ( .A(ram[2714]), .B(n12866), .Y(n2954) );
  OAI21X1 U5649 ( .A(n12710), .B(n12866), .C(n2955), .Y(n7152) );
  NAND2X1 U5650 ( .A(ram[2715]), .B(n12866), .Y(n2955) );
  OAI21X1 U5651 ( .A(n12704), .B(n12866), .C(n2956), .Y(n7153) );
  NAND2X1 U5652 ( .A(ram[2716]), .B(n12866), .Y(n2956) );
  OAI21X1 U5653 ( .A(n12698), .B(n12866), .C(n2957), .Y(n7154) );
  NAND2X1 U5654 ( .A(ram[2717]), .B(n12866), .Y(n2957) );
  OAI21X1 U5655 ( .A(n12695), .B(n12866), .C(n2958), .Y(n7155) );
  NAND2X1 U5656 ( .A(ram[2718]), .B(n12866), .Y(n2958) );
  OAI21X1 U5657 ( .A(n12689), .B(n12866), .C(n2959), .Y(n7156) );
  NAND2X1 U5658 ( .A(ram[2719]), .B(n12866), .Y(n2959) );
  OAI21X1 U5660 ( .A(n12778), .B(n12865), .C(n2961), .Y(n7157) );
  NAND2X1 U5661 ( .A(ram[2720]), .B(n12865), .Y(n2961) );
  OAI21X1 U5662 ( .A(n12772), .B(n12865), .C(n2962), .Y(n7158) );
  NAND2X1 U5663 ( .A(ram[2721]), .B(n12865), .Y(n2962) );
  OAI21X1 U5664 ( .A(n12762), .B(n12865), .C(n2963), .Y(n7159) );
  NAND2X1 U5665 ( .A(ram[2722]), .B(n12865), .Y(n2963) );
  OAI21X1 U5666 ( .A(n12756), .B(n12865), .C(n2964), .Y(n7160) );
  NAND2X1 U5667 ( .A(ram[2723]), .B(n12865), .Y(n2964) );
  OAI21X1 U5668 ( .A(n12750), .B(n12865), .C(n2965), .Y(n7161) );
  NAND2X1 U5669 ( .A(ram[2724]), .B(n12865), .Y(n2965) );
  OAI21X1 U5670 ( .A(n12744), .B(n12865), .C(n2966), .Y(n7162) );
  NAND2X1 U5671 ( .A(ram[2725]), .B(n12865), .Y(n2966) );
  OAI21X1 U5672 ( .A(n12738), .B(n12865), .C(n2967), .Y(n7163) );
  NAND2X1 U5673 ( .A(ram[2726]), .B(n12865), .Y(n2967) );
  OAI21X1 U5674 ( .A(n12732), .B(n12865), .C(n2968), .Y(n7164) );
  NAND2X1 U5675 ( .A(ram[2727]), .B(n12865), .Y(n2968) );
  OAI21X1 U5676 ( .A(n12726), .B(n12865), .C(n2969), .Y(n7165) );
  NAND2X1 U5677 ( .A(ram[2728]), .B(n12865), .Y(n2969) );
  OAI21X1 U5678 ( .A(n12720), .B(n12865), .C(n2970), .Y(n7166) );
  NAND2X1 U5679 ( .A(ram[2729]), .B(n12865), .Y(n2970) );
  OAI21X1 U5680 ( .A(n12714), .B(n12865), .C(n2971), .Y(n7167) );
  NAND2X1 U5681 ( .A(ram[2730]), .B(n12865), .Y(n2971) );
  OAI21X1 U5682 ( .A(n12708), .B(n12865), .C(n2972), .Y(n7168) );
  NAND2X1 U5683 ( .A(ram[2731]), .B(n12865), .Y(n2972) );
  OAI21X1 U5684 ( .A(n12702), .B(n12865), .C(n2973), .Y(n7169) );
  NAND2X1 U5685 ( .A(ram[2732]), .B(n12865), .Y(n2973) );
  OAI21X1 U5686 ( .A(n12696), .B(n12865), .C(n2974), .Y(n7170) );
  NAND2X1 U5687 ( .A(ram[2733]), .B(n12865), .Y(n2974) );
  OAI21X1 U5688 ( .A(n12694), .B(n12865), .C(n2975), .Y(n7171) );
  NAND2X1 U5689 ( .A(ram[2734]), .B(n12865), .Y(n2975) );
  OAI21X1 U5690 ( .A(n12688), .B(n12865), .C(n2976), .Y(n7172) );
  NAND2X1 U5691 ( .A(ram[2735]), .B(n12865), .Y(n2976) );
  OAI21X1 U5693 ( .A(n12777), .B(n12864), .C(n2978), .Y(n7173) );
  NAND2X1 U5694 ( .A(ram[2736]), .B(n12864), .Y(n2978) );
  OAI21X1 U5695 ( .A(n12771), .B(n12864), .C(n2979), .Y(n7174) );
  NAND2X1 U5696 ( .A(ram[2737]), .B(n12864), .Y(n2979) );
  OAI21X1 U5697 ( .A(n12763), .B(n12864), .C(n2980), .Y(n7175) );
  NAND2X1 U5698 ( .A(ram[2738]), .B(n12864), .Y(n2980) );
  OAI21X1 U5699 ( .A(n12757), .B(n12864), .C(n2981), .Y(n7176) );
  NAND2X1 U5700 ( .A(ram[2739]), .B(n12864), .Y(n2981) );
  OAI21X1 U5701 ( .A(n12751), .B(n12864), .C(n2982), .Y(n7177) );
  NAND2X1 U5702 ( .A(ram[2740]), .B(n12864), .Y(n2982) );
  OAI21X1 U5703 ( .A(n12745), .B(n12864), .C(n2983), .Y(n7178) );
  NAND2X1 U5704 ( .A(ram[2741]), .B(n12864), .Y(n2983) );
  OAI21X1 U5705 ( .A(n12739), .B(n12864), .C(n2984), .Y(n7179) );
  NAND2X1 U5706 ( .A(ram[2742]), .B(n12864), .Y(n2984) );
  OAI21X1 U5707 ( .A(n12733), .B(n12864), .C(n2985), .Y(n7180) );
  NAND2X1 U5708 ( .A(ram[2743]), .B(n12864), .Y(n2985) );
  OAI21X1 U5709 ( .A(n12727), .B(n12864), .C(n2986), .Y(n7181) );
  NAND2X1 U5710 ( .A(ram[2744]), .B(n12864), .Y(n2986) );
  OAI21X1 U5711 ( .A(n12721), .B(n12864), .C(n2987), .Y(n7182) );
  NAND2X1 U5712 ( .A(ram[2745]), .B(n12864), .Y(n2987) );
  OAI21X1 U5713 ( .A(n12715), .B(n12864), .C(n2988), .Y(n7183) );
  NAND2X1 U5714 ( .A(ram[2746]), .B(n12864), .Y(n2988) );
  OAI21X1 U5715 ( .A(n12709), .B(n12864), .C(n2989), .Y(n7184) );
  NAND2X1 U5716 ( .A(ram[2747]), .B(n12864), .Y(n2989) );
  OAI21X1 U5717 ( .A(n12703), .B(n12864), .C(n2990), .Y(n7185) );
  NAND2X1 U5718 ( .A(ram[2748]), .B(n12864), .Y(n2990) );
  OAI21X1 U5719 ( .A(n12697), .B(n12864), .C(n2991), .Y(n7186) );
  NAND2X1 U5720 ( .A(ram[2749]), .B(n12864), .Y(n2991) );
  OAI21X1 U5721 ( .A(n12693), .B(n12864), .C(n2992), .Y(n7187) );
  NAND2X1 U5722 ( .A(ram[2750]), .B(n12864), .Y(n2992) );
  OAI21X1 U5723 ( .A(n12687), .B(n12864), .C(n2993), .Y(n7188) );
  NAND2X1 U5724 ( .A(ram[2751]), .B(n12864), .Y(n2993) );
  OAI21X1 U5726 ( .A(n12775), .B(n12863), .C(n2995), .Y(n7189) );
  NAND2X1 U5727 ( .A(ram[2752]), .B(n12863), .Y(n2995) );
  OAI21X1 U5728 ( .A(n12769), .B(n12863), .C(n2996), .Y(n7190) );
  NAND2X1 U5729 ( .A(ram[2753]), .B(n12863), .Y(n2996) );
  OAI21X1 U5730 ( .A(n13069), .B(n12863), .C(n2997), .Y(n7191) );
  NAND2X1 U5731 ( .A(ram[2754]), .B(n12863), .Y(n2997) );
  OAI21X1 U5732 ( .A(n13068), .B(n12863), .C(n2998), .Y(n7192) );
  NAND2X1 U5733 ( .A(ram[2755]), .B(n12863), .Y(n2998) );
  OAI21X1 U5734 ( .A(n13067), .B(n12863), .C(n2999), .Y(n7193) );
  NAND2X1 U5735 ( .A(ram[2756]), .B(n12863), .Y(n2999) );
  OAI21X1 U5736 ( .A(n13066), .B(n12863), .C(n3000), .Y(n7194) );
  NAND2X1 U5737 ( .A(ram[2757]), .B(n12863), .Y(n3000) );
  OAI21X1 U5738 ( .A(n13065), .B(n12863), .C(n3001), .Y(n7195) );
  NAND2X1 U5739 ( .A(ram[2758]), .B(n12863), .Y(n3001) );
  OAI21X1 U5740 ( .A(n13064), .B(n12863), .C(n3002), .Y(n7196) );
  NAND2X1 U5741 ( .A(ram[2759]), .B(n12863), .Y(n3002) );
  OAI21X1 U5742 ( .A(n13063), .B(n12863), .C(n3003), .Y(n7197) );
  NAND2X1 U5743 ( .A(ram[2760]), .B(n12863), .Y(n3003) );
  OAI21X1 U5744 ( .A(n13062), .B(n12863), .C(n3004), .Y(n7198) );
  NAND2X1 U5745 ( .A(ram[2761]), .B(n12863), .Y(n3004) );
  OAI21X1 U5746 ( .A(n13061), .B(n12863), .C(n3005), .Y(n7199) );
  NAND2X1 U5747 ( .A(ram[2762]), .B(n12863), .Y(n3005) );
  OAI21X1 U5748 ( .A(n13060), .B(n12863), .C(n3006), .Y(n7200) );
  NAND2X1 U5749 ( .A(ram[2763]), .B(n12863), .Y(n3006) );
  OAI21X1 U5750 ( .A(n13059), .B(n12863), .C(n3007), .Y(n7201) );
  NAND2X1 U5751 ( .A(ram[2764]), .B(n12863), .Y(n3007) );
  OAI21X1 U5752 ( .A(n13058), .B(n12863), .C(n3008), .Y(n7202) );
  NAND2X1 U5753 ( .A(ram[2765]), .B(n12863), .Y(n3008) );
  OAI21X1 U5754 ( .A(n12691), .B(n12863), .C(n3009), .Y(n7203) );
  NAND2X1 U5755 ( .A(ram[2766]), .B(n12863), .Y(n3009) );
  OAI21X1 U5756 ( .A(n12685), .B(n12863), .C(n3010), .Y(n7204) );
  NAND2X1 U5757 ( .A(ram[2767]), .B(n12863), .Y(n3010) );
  OAI21X1 U5759 ( .A(n12777), .B(n12862), .C(n3012), .Y(n7205) );
  NAND2X1 U5760 ( .A(ram[2768]), .B(n12862), .Y(n3012) );
  OAI21X1 U5761 ( .A(n12771), .B(n12862), .C(n3013), .Y(n7206) );
  NAND2X1 U5762 ( .A(ram[2769]), .B(n12862), .Y(n3013) );
  OAI21X1 U5763 ( .A(n12762), .B(n12862), .C(n3014), .Y(n7207) );
  NAND2X1 U5764 ( .A(ram[2770]), .B(n12862), .Y(n3014) );
  OAI21X1 U5765 ( .A(n12756), .B(n12862), .C(n3015), .Y(n7208) );
  NAND2X1 U5766 ( .A(ram[2771]), .B(n12862), .Y(n3015) );
  OAI21X1 U5767 ( .A(n12750), .B(n12862), .C(n3016), .Y(n7209) );
  NAND2X1 U5768 ( .A(ram[2772]), .B(n12862), .Y(n3016) );
  OAI21X1 U5769 ( .A(n12744), .B(n12862), .C(n3017), .Y(n7210) );
  NAND2X1 U5770 ( .A(ram[2773]), .B(n12862), .Y(n3017) );
  OAI21X1 U5771 ( .A(n12738), .B(n12862), .C(n3018), .Y(n7211) );
  NAND2X1 U5772 ( .A(ram[2774]), .B(n12862), .Y(n3018) );
  OAI21X1 U5773 ( .A(n12732), .B(n12862), .C(n3019), .Y(n7212) );
  NAND2X1 U5774 ( .A(ram[2775]), .B(n12862), .Y(n3019) );
  OAI21X1 U5775 ( .A(n12726), .B(n12862), .C(n3020), .Y(n7213) );
  NAND2X1 U5776 ( .A(ram[2776]), .B(n12862), .Y(n3020) );
  OAI21X1 U5777 ( .A(n12720), .B(n12862), .C(n3021), .Y(n7214) );
  NAND2X1 U5778 ( .A(ram[2777]), .B(n12862), .Y(n3021) );
  OAI21X1 U5779 ( .A(n12714), .B(n12862), .C(n3022), .Y(n7215) );
  NAND2X1 U5780 ( .A(ram[2778]), .B(n12862), .Y(n3022) );
  OAI21X1 U5781 ( .A(n12708), .B(n12862), .C(n3023), .Y(n7216) );
  NAND2X1 U5782 ( .A(ram[2779]), .B(n12862), .Y(n3023) );
  OAI21X1 U5783 ( .A(n12702), .B(n12862), .C(n3024), .Y(n7217) );
  NAND2X1 U5784 ( .A(ram[2780]), .B(n12862), .Y(n3024) );
  OAI21X1 U5785 ( .A(n12696), .B(n12862), .C(n3025), .Y(n7218) );
  NAND2X1 U5786 ( .A(ram[2781]), .B(n12862), .Y(n3025) );
  OAI21X1 U5787 ( .A(n12693), .B(n12862), .C(n3026), .Y(n7219) );
  NAND2X1 U5788 ( .A(ram[2782]), .B(n12862), .Y(n3026) );
  OAI21X1 U5789 ( .A(n12687), .B(n12862), .C(n3027), .Y(n7220) );
  NAND2X1 U5790 ( .A(ram[2783]), .B(n12862), .Y(n3027) );
  OAI21X1 U5792 ( .A(n12775), .B(n12861), .C(n3029), .Y(n7221) );
  NAND2X1 U5793 ( .A(ram[2784]), .B(n12861), .Y(n3029) );
  OAI21X1 U5794 ( .A(n12769), .B(n12861), .C(n3030), .Y(n7222) );
  NAND2X1 U5795 ( .A(ram[2785]), .B(n12861), .Y(n3030) );
  OAI21X1 U5796 ( .A(n12762), .B(n12861), .C(n3031), .Y(n7223) );
  NAND2X1 U5797 ( .A(ram[2786]), .B(n12861), .Y(n3031) );
  OAI21X1 U5798 ( .A(n12756), .B(n12861), .C(n3032), .Y(n7224) );
  NAND2X1 U5799 ( .A(ram[2787]), .B(n12861), .Y(n3032) );
  OAI21X1 U5800 ( .A(n12750), .B(n12861), .C(n3033), .Y(n7225) );
  NAND2X1 U5801 ( .A(ram[2788]), .B(n12861), .Y(n3033) );
  OAI21X1 U5802 ( .A(n12744), .B(n12861), .C(n3034), .Y(n7226) );
  NAND2X1 U5803 ( .A(ram[2789]), .B(n12861), .Y(n3034) );
  OAI21X1 U5804 ( .A(n12738), .B(n12861), .C(n3035), .Y(n7227) );
  NAND2X1 U5805 ( .A(ram[2790]), .B(n12861), .Y(n3035) );
  OAI21X1 U5806 ( .A(n12732), .B(n12861), .C(n3036), .Y(n7228) );
  NAND2X1 U5807 ( .A(ram[2791]), .B(n12861), .Y(n3036) );
  OAI21X1 U5808 ( .A(n12726), .B(n12861), .C(n3037), .Y(n7229) );
  NAND2X1 U5809 ( .A(ram[2792]), .B(n12861), .Y(n3037) );
  OAI21X1 U5810 ( .A(n12720), .B(n12861), .C(n3038), .Y(n7230) );
  NAND2X1 U5811 ( .A(ram[2793]), .B(n12861), .Y(n3038) );
  OAI21X1 U5812 ( .A(n12714), .B(n12861), .C(n3039), .Y(n7231) );
  NAND2X1 U5813 ( .A(ram[2794]), .B(n12861), .Y(n3039) );
  OAI21X1 U5814 ( .A(n12708), .B(n12861), .C(n3040), .Y(n7232) );
  NAND2X1 U5815 ( .A(ram[2795]), .B(n12861), .Y(n3040) );
  OAI21X1 U5816 ( .A(n12702), .B(n12861), .C(n3041), .Y(n7233) );
  NAND2X1 U5817 ( .A(ram[2796]), .B(n12861), .Y(n3041) );
  OAI21X1 U5818 ( .A(n12696), .B(n12861), .C(n3042), .Y(n7234) );
  NAND2X1 U5819 ( .A(ram[2797]), .B(n12861), .Y(n3042) );
  OAI21X1 U5820 ( .A(n12691), .B(n12861), .C(n3043), .Y(n7235) );
  NAND2X1 U5821 ( .A(ram[2798]), .B(n12861), .Y(n3043) );
  OAI21X1 U5822 ( .A(n12685), .B(n12861), .C(n3044), .Y(n7236) );
  NAND2X1 U5823 ( .A(ram[2799]), .B(n12861), .Y(n3044) );
  OAI21X1 U5825 ( .A(n12778), .B(n12860), .C(n3046), .Y(n7237) );
  NAND2X1 U5826 ( .A(ram[2800]), .B(n12860), .Y(n3046) );
  OAI21X1 U5827 ( .A(n12772), .B(n12860), .C(n3047), .Y(n7238) );
  NAND2X1 U5828 ( .A(ram[2801]), .B(n12860), .Y(n3047) );
  OAI21X1 U5829 ( .A(n12763), .B(n12860), .C(n3048), .Y(n7239) );
  NAND2X1 U5830 ( .A(ram[2802]), .B(n12860), .Y(n3048) );
  OAI21X1 U5831 ( .A(n12757), .B(n12860), .C(n3049), .Y(n7240) );
  NAND2X1 U5832 ( .A(ram[2803]), .B(n12860), .Y(n3049) );
  OAI21X1 U5833 ( .A(n12751), .B(n12860), .C(n3050), .Y(n7241) );
  NAND2X1 U5834 ( .A(ram[2804]), .B(n12860), .Y(n3050) );
  OAI21X1 U5835 ( .A(n12745), .B(n12860), .C(n3051), .Y(n7242) );
  NAND2X1 U5836 ( .A(ram[2805]), .B(n12860), .Y(n3051) );
  OAI21X1 U5837 ( .A(n12739), .B(n12860), .C(n3052), .Y(n7243) );
  NAND2X1 U5838 ( .A(ram[2806]), .B(n12860), .Y(n3052) );
  OAI21X1 U5839 ( .A(n12733), .B(n12860), .C(n3053), .Y(n7244) );
  NAND2X1 U5840 ( .A(ram[2807]), .B(n12860), .Y(n3053) );
  OAI21X1 U5841 ( .A(n12727), .B(n12860), .C(n3054), .Y(n7245) );
  NAND2X1 U5842 ( .A(ram[2808]), .B(n12860), .Y(n3054) );
  OAI21X1 U5843 ( .A(n12721), .B(n12860), .C(n3055), .Y(n7246) );
  NAND2X1 U5844 ( .A(ram[2809]), .B(n12860), .Y(n3055) );
  OAI21X1 U5845 ( .A(n12715), .B(n12860), .C(n3056), .Y(n7247) );
  NAND2X1 U5846 ( .A(ram[2810]), .B(n12860), .Y(n3056) );
  OAI21X1 U5847 ( .A(n12709), .B(n12860), .C(n3057), .Y(n7248) );
  NAND2X1 U5848 ( .A(ram[2811]), .B(n12860), .Y(n3057) );
  OAI21X1 U5849 ( .A(n12703), .B(n12860), .C(n3058), .Y(n7249) );
  NAND2X1 U5850 ( .A(ram[2812]), .B(n12860), .Y(n3058) );
  OAI21X1 U5851 ( .A(n12697), .B(n12860), .C(n3059), .Y(n7250) );
  NAND2X1 U5852 ( .A(ram[2813]), .B(n12860), .Y(n3059) );
  OAI21X1 U5853 ( .A(n12694), .B(n12860), .C(n3060), .Y(n7251) );
  NAND2X1 U5854 ( .A(ram[2814]), .B(n12860), .Y(n3060) );
  OAI21X1 U5855 ( .A(n12688), .B(n12860), .C(n3061), .Y(n7252) );
  NAND2X1 U5856 ( .A(ram[2815]), .B(n12860), .Y(n3061) );
  NAND3X1 U5858 ( .A(n875), .B(mem_write_en), .C(n2516), .Y(n3062) );
  OAI21X1 U5859 ( .A(n12774), .B(n12859), .C(n3064), .Y(n7253) );
  NAND2X1 U5860 ( .A(ram[2816]), .B(n12859), .Y(n3064) );
  OAI21X1 U5861 ( .A(n12768), .B(n12859), .C(n3065), .Y(n7254) );
  NAND2X1 U5862 ( .A(ram[2817]), .B(n12859), .Y(n3065) );
  OAI21X1 U5863 ( .A(n12763), .B(n12859), .C(n3066), .Y(n7255) );
  NAND2X1 U5864 ( .A(ram[2818]), .B(n12859), .Y(n3066) );
  OAI21X1 U5865 ( .A(n12757), .B(n12859), .C(n3067), .Y(n7256) );
  NAND2X1 U5866 ( .A(ram[2819]), .B(n12859), .Y(n3067) );
  OAI21X1 U5867 ( .A(n12751), .B(n12859), .C(n3068), .Y(n7257) );
  NAND2X1 U5868 ( .A(ram[2820]), .B(n12859), .Y(n3068) );
  OAI21X1 U5869 ( .A(n12745), .B(n12859), .C(n3069), .Y(n7258) );
  NAND2X1 U5870 ( .A(ram[2821]), .B(n12859), .Y(n3069) );
  OAI21X1 U5871 ( .A(n12739), .B(n12859), .C(n3070), .Y(n7259) );
  NAND2X1 U5872 ( .A(ram[2822]), .B(n12859), .Y(n3070) );
  OAI21X1 U5873 ( .A(n12733), .B(n12859), .C(n3071), .Y(n7260) );
  NAND2X1 U5874 ( .A(ram[2823]), .B(n12859), .Y(n3071) );
  OAI21X1 U5875 ( .A(n12727), .B(n12859), .C(n3072), .Y(n7261) );
  NAND2X1 U5876 ( .A(ram[2824]), .B(n12859), .Y(n3072) );
  OAI21X1 U5877 ( .A(n12721), .B(n12859), .C(n3073), .Y(n7262) );
  NAND2X1 U5878 ( .A(ram[2825]), .B(n12859), .Y(n3073) );
  OAI21X1 U5879 ( .A(n12715), .B(n12859), .C(n3074), .Y(n7263) );
  NAND2X1 U5880 ( .A(ram[2826]), .B(n12859), .Y(n3074) );
  OAI21X1 U5881 ( .A(n12709), .B(n12859), .C(n3075), .Y(n7264) );
  NAND2X1 U5882 ( .A(ram[2827]), .B(n12859), .Y(n3075) );
  OAI21X1 U5883 ( .A(n12703), .B(n12859), .C(n3076), .Y(n7265) );
  NAND2X1 U5884 ( .A(ram[2828]), .B(n12859), .Y(n3076) );
  OAI21X1 U5885 ( .A(n12697), .B(n12859), .C(n3077), .Y(n7266) );
  NAND2X1 U5886 ( .A(ram[2829]), .B(n12859), .Y(n3077) );
  OAI21X1 U5887 ( .A(n12690), .B(n12859), .C(n3078), .Y(n7267) );
  NAND2X1 U5888 ( .A(ram[2830]), .B(n12859), .Y(n3078) );
  OAI21X1 U5889 ( .A(n12684), .B(n12859), .C(n3079), .Y(n7268) );
  NAND2X1 U5890 ( .A(ram[2831]), .B(n12859), .Y(n3079) );
  OAI21X1 U5892 ( .A(n12774), .B(n12858), .C(n3081), .Y(n7269) );
  NAND2X1 U5893 ( .A(ram[2832]), .B(n12858), .Y(n3081) );
  OAI21X1 U5894 ( .A(n12768), .B(n12858), .C(n3082), .Y(n7270) );
  NAND2X1 U5895 ( .A(ram[2833]), .B(n12858), .Y(n3082) );
  OAI21X1 U5896 ( .A(n12763), .B(n12858), .C(n3083), .Y(n7271) );
  NAND2X1 U5897 ( .A(ram[2834]), .B(n12858), .Y(n3083) );
  OAI21X1 U5898 ( .A(n12757), .B(n12858), .C(n3084), .Y(n7272) );
  NAND2X1 U5899 ( .A(ram[2835]), .B(n12858), .Y(n3084) );
  OAI21X1 U5900 ( .A(n12751), .B(n12858), .C(n3085), .Y(n7273) );
  NAND2X1 U5901 ( .A(ram[2836]), .B(n12858), .Y(n3085) );
  OAI21X1 U5902 ( .A(n12745), .B(n12858), .C(n3086), .Y(n7274) );
  NAND2X1 U5903 ( .A(ram[2837]), .B(n12858), .Y(n3086) );
  OAI21X1 U5904 ( .A(n12739), .B(n12858), .C(n3087), .Y(n7275) );
  NAND2X1 U5905 ( .A(ram[2838]), .B(n12858), .Y(n3087) );
  OAI21X1 U5906 ( .A(n12733), .B(n12858), .C(n3088), .Y(n7276) );
  NAND2X1 U5907 ( .A(ram[2839]), .B(n12858), .Y(n3088) );
  OAI21X1 U5908 ( .A(n12727), .B(n12858), .C(n3089), .Y(n7277) );
  NAND2X1 U5909 ( .A(ram[2840]), .B(n12858), .Y(n3089) );
  OAI21X1 U5910 ( .A(n12721), .B(n12858), .C(n3090), .Y(n7278) );
  NAND2X1 U5911 ( .A(ram[2841]), .B(n12858), .Y(n3090) );
  OAI21X1 U5912 ( .A(n12715), .B(n12858), .C(n3091), .Y(n7279) );
  NAND2X1 U5913 ( .A(ram[2842]), .B(n12858), .Y(n3091) );
  OAI21X1 U5914 ( .A(n12709), .B(n12858), .C(n3092), .Y(n7280) );
  NAND2X1 U5915 ( .A(ram[2843]), .B(n12858), .Y(n3092) );
  OAI21X1 U5916 ( .A(n12703), .B(n12858), .C(n3093), .Y(n7281) );
  NAND2X1 U5917 ( .A(ram[2844]), .B(n12858), .Y(n3093) );
  OAI21X1 U5918 ( .A(n12697), .B(n12858), .C(n3094), .Y(n7282) );
  NAND2X1 U5919 ( .A(ram[2845]), .B(n12858), .Y(n3094) );
  OAI21X1 U5920 ( .A(n12690), .B(n12858), .C(n3095), .Y(n7283) );
  NAND2X1 U5921 ( .A(ram[2846]), .B(n12858), .Y(n3095) );
  OAI21X1 U5922 ( .A(n12684), .B(n12858), .C(n3096), .Y(n7284) );
  NAND2X1 U5923 ( .A(ram[2847]), .B(n12858), .Y(n3096) );
  OAI21X1 U5925 ( .A(n12775), .B(n12857), .C(n3098), .Y(n7285) );
  NAND2X1 U5926 ( .A(ram[2848]), .B(n12857), .Y(n3098) );
  OAI21X1 U5927 ( .A(n12769), .B(n12857), .C(n3099), .Y(n7286) );
  NAND2X1 U5928 ( .A(ram[2849]), .B(n12857), .Y(n3099) );
  OAI21X1 U5929 ( .A(n12762), .B(n12857), .C(n3100), .Y(n7287) );
  NAND2X1 U5930 ( .A(ram[2850]), .B(n12857), .Y(n3100) );
  OAI21X1 U5931 ( .A(n12756), .B(n12857), .C(n3101), .Y(n7288) );
  NAND2X1 U5932 ( .A(ram[2851]), .B(n12857), .Y(n3101) );
  OAI21X1 U5933 ( .A(n12750), .B(n12857), .C(n3102), .Y(n7289) );
  NAND2X1 U5934 ( .A(ram[2852]), .B(n12857), .Y(n3102) );
  OAI21X1 U5935 ( .A(n12744), .B(n12857), .C(n3103), .Y(n7290) );
  NAND2X1 U5936 ( .A(ram[2853]), .B(n12857), .Y(n3103) );
  OAI21X1 U5937 ( .A(n12738), .B(n12857), .C(n3104), .Y(n7291) );
  NAND2X1 U5938 ( .A(ram[2854]), .B(n12857), .Y(n3104) );
  OAI21X1 U5939 ( .A(n12732), .B(n12857), .C(n3105), .Y(n7292) );
  NAND2X1 U5940 ( .A(ram[2855]), .B(n12857), .Y(n3105) );
  OAI21X1 U5941 ( .A(n12726), .B(n12857), .C(n3106), .Y(n7293) );
  NAND2X1 U5942 ( .A(ram[2856]), .B(n12857), .Y(n3106) );
  OAI21X1 U5943 ( .A(n12720), .B(n12857), .C(n3107), .Y(n7294) );
  NAND2X1 U5944 ( .A(ram[2857]), .B(n12857), .Y(n3107) );
  OAI21X1 U5945 ( .A(n12714), .B(n12857), .C(n3108), .Y(n7295) );
  NAND2X1 U5946 ( .A(ram[2858]), .B(n12857), .Y(n3108) );
  OAI21X1 U5947 ( .A(n12708), .B(n12857), .C(n3109), .Y(n7296) );
  NAND2X1 U5948 ( .A(ram[2859]), .B(n12857), .Y(n3109) );
  OAI21X1 U5949 ( .A(n12702), .B(n12857), .C(n3110), .Y(n7297) );
  NAND2X1 U5950 ( .A(ram[2860]), .B(n12857), .Y(n3110) );
  OAI21X1 U5951 ( .A(n12696), .B(n12857), .C(n3111), .Y(n7298) );
  NAND2X1 U5952 ( .A(ram[2861]), .B(n12857), .Y(n3111) );
  OAI21X1 U5953 ( .A(n12691), .B(n12857), .C(n3112), .Y(n7299) );
  NAND2X1 U5954 ( .A(ram[2862]), .B(n12857), .Y(n3112) );
  OAI21X1 U5955 ( .A(n12685), .B(n12857), .C(n3113), .Y(n7300) );
  NAND2X1 U5956 ( .A(ram[2863]), .B(n12857), .Y(n3113) );
  OAI21X1 U5958 ( .A(n13071), .B(n12856), .C(n3115), .Y(n7301) );
  NAND2X1 U5959 ( .A(ram[2864]), .B(n12856), .Y(n3115) );
  OAI21X1 U5960 ( .A(n13070), .B(n12856), .C(n3116), .Y(n7302) );
  NAND2X1 U5961 ( .A(ram[2865]), .B(n12856), .Y(n3116) );
  OAI21X1 U5962 ( .A(n12763), .B(n12856), .C(n3117), .Y(n7303) );
  NAND2X1 U5963 ( .A(ram[2866]), .B(n12856), .Y(n3117) );
  OAI21X1 U5964 ( .A(n12757), .B(n12856), .C(n3118), .Y(n7304) );
  NAND2X1 U5965 ( .A(ram[2867]), .B(n12856), .Y(n3118) );
  OAI21X1 U5966 ( .A(n12751), .B(n12856), .C(n3119), .Y(n7305) );
  NAND2X1 U5967 ( .A(ram[2868]), .B(n12856), .Y(n3119) );
  OAI21X1 U5968 ( .A(n12745), .B(n12856), .C(n3120), .Y(n7306) );
  NAND2X1 U5969 ( .A(ram[2869]), .B(n12856), .Y(n3120) );
  OAI21X1 U5970 ( .A(n12739), .B(n12856), .C(n3121), .Y(n7307) );
  NAND2X1 U5971 ( .A(ram[2870]), .B(n12856), .Y(n3121) );
  OAI21X1 U5972 ( .A(n12733), .B(n12856), .C(n3122), .Y(n7308) );
  NAND2X1 U5973 ( .A(ram[2871]), .B(n12856), .Y(n3122) );
  OAI21X1 U5974 ( .A(n12727), .B(n12856), .C(n3123), .Y(n7309) );
  NAND2X1 U5975 ( .A(ram[2872]), .B(n12856), .Y(n3123) );
  OAI21X1 U5976 ( .A(n12721), .B(n12856), .C(n3124), .Y(n7310) );
  NAND2X1 U5977 ( .A(ram[2873]), .B(n12856), .Y(n3124) );
  OAI21X1 U5978 ( .A(n12715), .B(n12856), .C(n3125), .Y(n7311) );
  NAND2X1 U5979 ( .A(ram[2874]), .B(n12856), .Y(n3125) );
  OAI21X1 U5980 ( .A(n12709), .B(n12856), .C(n3126), .Y(n7312) );
  NAND2X1 U5981 ( .A(ram[2875]), .B(n12856), .Y(n3126) );
  OAI21X1 U5982 ( .A(n12703), .B(n12856), .C(n3127), .Y(n7313) );
  NAND2X1 U5983 ( .A(ram[2876]), .B(n12856), .Y(n3127) );
  OAI21X1 U5984 ( .A(n12697), .B(n12856), .C(n3128), .Y(n7314) );
  NAND2X1 U5985 ( .A(ram[2877]), .B(n12856), .Y(n3128) );
  OAI21X1 U5986 ( .A(n13057), .B(n12856), .C(n3129), .Y(n7315) );
  NAND2X1 U5987 ( .A(ram[2878]), .B(n12856), .Y(n3129) );
  OAI21X1 U5988 ( .A(n13056), .B(n12856), .C(n3130), .Y(n7316) );
  NAND2X1 U5989 ( .A(ram[2879]), .B(n12856), .Y(n3130) );
  OAI21X1 U5991 ( .A(n12777), .B(n12855), .C(n3132), .Y(n7317) );
  NAND2X1 U5992 ( .A(ram[2880]), .B(n12855), .Y(n3132) );
  OAI21X1 U5993 ( .A(n12771), .B(n12855), .C(n3133), .Y(n7318) );
  NAND2X1 U5994 ( .A(ram[2881]), .B(n12855), .Y(n3133) );
  OAI21X1 U5995 ( .A(n12762), .B(n12855), .C(n3134), .Y(n7319) );
  NAND2X1 U5996 ( .A(ram[2882]), .B(n12855), .Y(n3134) );
  OAI21X1 U5997 ( .A(n12756), .B(n12855), .C(n3135), .Y(n7320) );
  NAND2X1 U5998 ( .A(ram[2883]), .B(n12855), .Y(n3135) );
  OAI21X1 U5999 ( .A(n12750), .B(n12855), .C(n3136), .Y(n7321) );
  NAND2X1 U6000 ( .A(ram[2884]), .B(n12855), .Y(n3136) );
  OAI21X1 U6001 ( .A(n12744), .B(n12855), .C(n3137), .Y(n7322) );
  NAND2X1 U6002 ( .A(ram[2885]), .B(n12855), .Y(n3137) );
  OAI21X1 U6003 ( .A(n12738), .B(n12855), .C(n3138), .Y(n7323) );
  NAND2X1 U6004 ( .A(ram[2886]), .B(n12855), .Y(n3138) );
  OAI21X1 U6005 ( .A(n12732), .B(n12855), .C(n3139), .Y(n7324) );
  NAND2X1 U6006 ( .A(ram[2887]), .B(n12855), .Y(n3139) );
  OAI21X1 U6007 ( .A(n12726), .B(n12855), .C(n3140), .Y(n7325) );
  NAND2X1 U6008 ( .A(ram[2888]), .B(n12855), .Y(n3140) );
  OAI21X1 U6009 ( .A(n12720), .B(n12855), .C(n3141), .Y(n7326) );
  NAND2X1 U6010 ( .A(ram[2889]), .B(n12855), .Y(n3141) );
  OAI21X1 U6011 ( .A(n12714), .B(n12855), .C(n3142), .Y(n7327) );
  NAND2X1 U6012 ( .A(ram[2890]), .B(n12855), .Y(n3142) );
  OAI21X1 U6013 ( .A(n12708), .B(n12855), .C(n3143), .Y(n7328) );
  NAND2X1 U6014 ( .A(ram[2891]), .B(n12855), .Y(n3143) );
  OAI21X1 U6015 ( .A(n12702), .B(n12855), .C(n3144), .Y(n7329) );
  NAND2X1 U6016 ( .A(ram[2892]), .B(n12855), .Y(n3144) );
  OAI21X1 U6017 ( .A(n12696), .B(n12855), .C(n3145), .Y(n7330) );
  NAND2X1 U6018 ( .A(ram[2893]), .B(n12855), .Y(n3145) );
  OAI21X1 U6019 ( .A(n12693), .B(n12855), .C(n3146), .Y(n7331) );
  NAND2X1 U6020 ( .A(ram[2894]), .B(n12855), .Y(n3146) );
  OAI21X1 U6021 ( .A(n12687), .B(n12855), .C(n3147), .Y(n7332) );
  NAND2X1 U6022 ( .A(ram[2895]), .B(n12855), .Y(n3147) );
  OAI21X1 U6024 ( .A(n12776), .B(n12854), .C(n3149), .Y(n7333) );
  NAND2X1 U6025 ( .A(ram[2896]), .B(n12854), .Y(n3149) );
  OAI21X1 U6026 ( .A(n12770), .B(n12854), .C(n3150), .Y(n7334) );
  NAND2X1 U6027 ( .A(ram[2897]), .B(n12854), .Y(n3150) );
  OAI21X1 U6028 ( .A(n12766), .B(n12854), .C(n3151), .Y(n7335) );
  NAND2X1 U6029 ( .A(ram[2898]), .B(n12854), .Y(n3151) );
  OAI21X1 U6030 ( .A(n12760), .B(n12854), .C(n3152), .Y(n7336) );
  NAND2X1 U6031 ( .A(ram[2899]), .B(n12854), .Y(n3152) );
  OAI21X1 U6032 ( .A(n12754), .B(n12854), .C(n3153), .Y(n7337) );
  NAND2X1 U6033 ( .A(ram[2900]), .B(n12854), .Y(n3153) );
  OAI21X1 U6034 ( .A(n12748), .B(n12854), .C(n3154), .Y(n7338) );
  NAND2X1 U6035 ( .A(ram[2901]), .B(n12854), .Y(n3154) );
  OAI21X1 U6036 ( .A(n12742), .B(n12854), .C(n3155), .Y(n7339) );
  NAND2X1 U6037 ( .A(ram[2902]), .B(n12854), .Y(n3155) );
  OAI21X1 U6038 ( .A(n12736), .B(n12854), .C(n3156), .Y(n7340) );
  NAND2X1 U6039 ( .A(ram[2903]), .B(n12854), .Y(n3156) );
  OAI21X1 U6040 ( .A(n12730), .B(n12854), .C(n3157), .Y(n7341) );
  NAND2X1 U6041 ( .A(ram[2904]), .B(n12854), .Y(n3157) );
  OAI21X1 U6042 ( .A(n12724), .B(n12854), .C(n3158), .Y(n7342) );
  NAND2X1 U6043 ( .A(ram[2905]), .B(n12854), .Y(n3158) );
  OAI21X1 U6044 ( .A(n12718), .B(n12854), .C(n3159), .Y(n7343) );
  NAND2X1 U6045 ( .A(ram[2906]), .B(n12854), .Y(n3159) );
  OAI21X1 U6046 ( .A(n12712), .B(n12854), .C(n3160), .Y(n7344) );
  NAND2X1 U6047 ( .A(ram[2907]), .B(n12854), .Y(n3160) );
  OAI21X1 U6048 ( .A(n12706), .B(n12854), .C(n3161), .Y(n7345) );
  NAND2X1 U6049 ( .A(ram[2908]), .B(n12854), .Y(n3161) );
  OAI21X1 U6050 ( .A(n12700), .B(n12854), .C(n3162), .Y(n7346) );
  NAND2X1 U6051 ( .A(ram[2909]), .B(n12854), .Y(n3162) );
  OAI21X1 U6052 ( .A(n12692), .B(n12854), .C(n3163), .Y(n7347) );
  NAND2X1 U6053 ( .A(ram[2910]), .B(n12854), .Y(n3163) );
  OAI21X1 U6054 ( .A(n12686), .B(n12854), .C(n3164), .Y(n7348) );
  NAND2X1 U6055 ( .A(ram[2911]), .B(n12854), .Y(n3164) );
  OAI21X1 U6057 ( .A(n12776), .B(n12853), .C(n3166), .Y(n7349) );
  NAND2X1 U6058 ( .A(ram[2912]), .B(n12853), .Y(n3166) );
  OAI21X1 U6059 ( .A(n12770), .B(n12853), .C(n3167), .Y(n7350) );
  NAND2X1 U6060 ( .A(ram[2913]), .B(n12853), .Y(n3167) );
  OAI21X1 U6061 ( .A(n12764), .B(n12853), .C(n3168), .Y(n7351) );
  NAND2X1 U6062 ( .A(ram[2914]), .B(n12853), .Y(n3168) );
  OAI21X1 U6063 ( .A(n12758), .B(n12853), .C(n3169), .Y(n7352) );
  NAND2X1 U6064 ( .A(ram[2915]), .B(n12853), .Y(n3169) );
  OAI21X1 U6065 ( .A(n12752), .B(n12853), .C(n3170), .Y(n7353) );
  NAND2X1 U6066 ( .A(ram[2916]), .B(n12853), .Y(n3170) );
  OAI21X1 U6067 ( .A(n12746), .B(n12853), .C(n3171), .Y(n7354) );
  NAND2X1 U6068 ( .A(ram[2917]), .B(n12853), .Y(n3171) );
  OAI21X1 U6069 ( .A(n12740), .B(n12853), .C(n3172), .Y(n7355) );
  NAND2X1 U6070 ( .A(ram[2918]), .B(n12853), .Y(n3172) );
  OAI21X1 U6071 ( .A(n12734), .B(n12853), .C(n3173), .Y(n7356) );
  NAND2X1 U6072 ( .A(ram[2919]), .B(n12853), .Y(n3173) );
  OAI21X1 U6073 ( .A(n12728), .B(n12853), .C(n3174), .Y(n7357) );
  NAND2X1 U6074 ( .A(ram[2920]), .B(n12853), .Y(n3174) );
  OAI21X1 U6075 ( .A(n12722), .B(n12853), .C(n3175), .Y(n7358) );
  NAND2X1 U6076 ( .A(ram[2921]), .B(n12853), .Y(n3175) );
  OAI21X1 U6077 ( .A(n12716), .B(n12853), .C(n3176), .Y(n7359) );
  NAND2X1 U6078 ( .A(ram[2922]), .B(n12853), .Y(n3176) );
  OAI21X1 U6079 ( .A(n12710), .B(n12853), .C(n3177), .Y(n7360) );
  NAND2X1 U6080 ( .A(ram[2923]), .B(n12853), .Y(n3177) );
  OAI21X1 U6081 ( .A(n12704), .B(n12853), .C(n3178), .Y(n7361) );
  NAND2X1 U6082 ( .A(ram[2924]), .B(n12853), .Y(n3178) );
  OAI21X1 U6083 ( .A(n12698), .B(n12853), .C(n3179), .Y(n7362) );
  NAND2X1 U6084 ( .A(ram[2925]), .B(n12853), .Y(n3179) );
  OAI21X1 U6085 ( .A(n12692), .B(n12853), .C(n3180), .Y(n7363) );
  NAND2X1 U6086 ( .A(ram[2926]), .B(n12853), .Y(n3180) );
  OAI21X1 U6087 ( .A(n12686), .B(n12853), .C(n3181), .Y(n7364) );
  NAND2X1 U6088 ( .A(ram[2927]), .B(n12853), .Y(n3181) );
  OAI21X1 U6090 ( .A(n12776), .B(n12852), .C(n3183), .Y(n7365) );
  NAND2X1 U6091 ( .A(ram[2928]), .B(n12852), .Y(n3183) );
  OAI21X1 U6092 ( .A(n12770), .B(n12852), .C(n3184), .Y(n7366) );
  NAND2X1 U6093 ( .A(ram[2929]), .B(n12852), .Y(n3184) );
  OAI21X1 U6094 ( .A(n12764), .B(n12852), .C(n3185), .Y(n7367) );
  NAND2X1 U6095 ( .A(ram[2930]), .B(n12852), .Y(n3185) );
  OAI21X1 U6096 ( .A(n12758), .B(n12852), .C(n3186), .Y(n7368) );
  NAND2X1 U6097 ( .A(ram[2931]), .B(n12852), .Y(n3186) );
  OAI21X1 U6098 ( .A(n12752), .B(n12852), .C(n3187), .Y(n7369) );
  NAND2X1 U6099 ( .A(ram[2932]), .B(n12852), .Y(n3187) );
  OAI21X1 U6100 ( .A(n12746), .B(n12852), .C(n3188), .Y(n7370) );
  NAND2X1 U6101 ( .A(ram[2933]), .B(n12852), .Y(n3188) );
  OAI21X1 U6102 ( .A(n12740), .B(n12852), .C(n3189), .Y(n7371) );
  NAND2X1 U6103 ( .A(ram[2934]), .B(n12852), .Y(n3189) );
  OAI21X1 U6104 ( .A(n12734), .B(n12852), .C(n3190), .Y(n7372) );
  NAND2X1 U6105 ( .A(ram[2935]), .B(n12852), .Y(n3190) );
  OAI21X1 U6106 ( .A(n12728), .B(n12852), .C(n3191), .Y(n7373) );
  NAND2X1 U6107 ( .A(ram[2936]), .B(n12852), .Y(n3191) );
  OAI21X1 U6108 ( .A(n12722), .B(n12852), .C(n3192), .Y(n7374) );
  NAND2X1 U6109 ( .A(ram[2937]), .B(n12852), .Y(n3192) );
  OAI21X1 U6110 ( .A(n12716), .B(n12852), .C(n3193), .Y(n7375) );
  NAND2X1 U6111 ( .A(ram[2938]), .B(n12852), .Y(n3193) );
  OAI21X1 U6112 ( .A(n12710), .B(n12852), .C(n3194), .Y(n7376) );
  NAND2X1 U6113 ( .A(ram[2939]), .B(n12852), .Y(n3194) );
  OAI21X1 U6114 ( .A(n12704), .B(n12852), .C(n3195), .Y(n7377) );
  NAND2X1 U6115 ( .A(ram[2940]), .B(n12852), .Y(n3195) );
  OAI21X1 U6116 ( .A(n12698), .B(n12852), .C(n3196), .Y(n7378) );
  NAND2X1 U6117 ( .A(ram[2941]), .B(n12852), .Y(n3196) );
  OAI21X1 U6118 ( .A(n12692), .B(n12852), .C(n3197), .Y(n7379) );
  NAND2X1 U6119 ( .A(ram[2942]), .B(n12852), .Y(n3197) );
  OAI21X1 U6120 ( .A(n12686), .B(n12852), .C(n3198), .Y(n7380) );
  NAND2X1 U6121 ( .A(ram[2943]), .B(n12852), .Y(n3198) );
  OAI21X1 U6123 ( .A(n12776), .B(n12851), .C(n3200), .Y(n7381) );
  NAND2X1 U6124 ( .A(ram[2944]), .B(n12851), .Y(n3200) );
  OAI21X1 U6125 ( .A(n12770), .B(n12851), .C(n3201), .Y(n7382) );
  NAND2X1 U6126 ( .A(ram[2945]), .B(n12851), .Y(n3201) );
  OAI21X1 U6127 ( .A(n12764), .B(n12851), .C(n3202), .Y(n7383) );
  NAND2X1 U6128 ( .A(ram[2946]), .B(n12851), .Y(n3202) );
  OAI21X1 U6129 ( .A(n12758), .B(n12851), .C(n3203), .Y(n7384) );
  NAND2X1 U6130 ( .A(ram[2947]), .B(n12851), .Y(n3203) );
  OAI21X1 U6131 ( .A(n12752), .B(n12851), .C(n3204), .Y(n7385) );
  NAND2X1 U6132 ( .A(ram[2948]), .B(n12851), .Y(n3204) );
  OAI21X1 U6133 ( .A(n12746), .B(n12851), .C(n3205), .Y(n7386) );
  NAND2X1 U6134 ( .A(ram[2949]), .B(n12851), .Y(n3205) );
  OAI21X1 U6135 ( .A(n12740), .B(n12851), .C(n3206), .Y(n7387) );
  NAND2X1 U6136 ( .A(ram[2950]), .B(n12851), .Y(n3206) );
  OAI21X1 U6137 ( .A(n12734), .B(n12851), .C(n3207), .Y(n7388) );
  NAND2X1 U6138 ( .A(ram[2951]), .B(n12851), .Y(n3207) );
  OAI21X1 U6139 ( .A(n12728), .B(n12851), .C(n3208), .Y(n7389) );
  NAND2X1 U6140 ( .A(ram[2952]), .B(n12851), .Y(n3208) );
  OAI21X1 U6141 ( .A(n12722), .B(n12851), .C(n3209), .Y(n7390) );
  NAND2X1 U6142 ( .A(ram[2953]), .B(n12851), .Y(n3209) );
  OAI21X1 U6143 ( .A(n12716), .B(n12851), .C(n3210), .Y(n7391) );
  NAND2X1 U6144 ( .A(ram[2954]), .B(n12851), .Y(n3210) );
  OAI21X1 U6145 ( .A(n12710), .B(n12851), .C(n3211), .Y(n7392) );
  NAND2X1 U6146 ( .A(ram[2955]), .B(n12851), .Y(n3211) );
  OAI21X1 U6147 ( .A(n12704), .B(n12851), .C(n3212), .Y(n7393) );
  NAND2X1 U6148 ( .A(ram[2956]), .B(n12851), .Y(n3212) );
  OAI21X1 U6149 ( .A(n12698), .B(n12851), .C(n3213), .Y(n7394) );
  NAND2X1 U6150 ( .A(ram[2957]), .B(n12851), .Y(n3213) );
  OAI21X1 U6151 ( .A(n12692), .B(n12851), .C(n3214), .Y(n7395) );
  NAND2X1 U6152 ( .A(ram[2958]), .B(n12851), .Y(n3214) );
  OAI21X1 U6153 ( .A(n12686), .B(n12851), .C(n3215), .Y(n7396) );
  NAND2X1 U6154 ( .A(ram[2959]), .B(n12851), .Y(n3215) );
  OAI21X1 U6156 ( .A(n12776), .B(n12850), .C(n3217), .Y(n7397) );
  NAND2X1 U6157 ( .A(ram[2960]), .B(n12850), .Y(n3217) );
  OAI21X1 U6158 ( .A(n12770), .B(n12850), .C(n3218), .Y(n7398) );
  NAND2X1 U6159 ( .A(ram[2961]), .B(n12850), .Y(n3218) );
  OAI21X1 U6160 ( .A(n12764), .B(n12850), .C(n3219), .Y(n7399) );
  NAND2X1 U6161 ( .A(ram[2962]), .B(n12850), .Y(n3219) );
  OAI21X1 U6162 ( .A(n12758), .B(n12850), .C(n3220), .Y(n7400) );
  NAND2X1 U6163 ( .A(ram[2963]), .B(n12850), .Y(n3220) );
  OAI21X1 U6164 ( .A(n12752), .B(n12850), .C(n3221), .Y(n7401) );
  NAND2X1 U6165 ( .A(ram[2964]), .B(n12850), .Y(n3221) );
  OAI21X1 U6166 ( .A(n12746), .B(n12850), .C(n3222), .Y(n7402) );
  NAND2X1 U6167 ( .A(ram[2965]), .B(n12850), .Y(n3222) );
  OAI21X1 U6168 ( .A(n12740), .B(n12850), .C(n3223), .Y(n7403) );
  NAND2X1 U6169 ( .A(ram[2966]), .B(n12850), .Y(n3223) );
  OAI21X1 U6170 ( .A(n12734), .B(n12850), .C(n3224), .Y(n7404) );
  NAND2X1 U6171 ( .A(ram[2967]), .B(n12850), .Y(n3224) );
  OAI21X1 U6172 ( .A(n12728), .B(n12850), .C(n3225), .Y(n7405) );
  NAND2X1 U6173 ( .A(ram[2968]), .B(n12850), .Y(n3225) );
  OAI21X1 U6174 ( .A(n12722), .B(n12850), .C(n3226), .Y(n7406) );
  NAND2X1 U6175 ( .A(ram[2969]), .B(n12850), .Y(n3226) );
  OAI21X1 U6176 ( .A(n12716), .B(n12850), .C(n3227), .Y(n7407) );
  NAND2X1 U6177 ( .A(ram[2970]), .B(n12850), .Y(n3227) );
  OAI21X1 U6178 ( .A(n12710), .B(n12850), .C(n3228), .Y(n7408) );
  NAND2X1 U6179 ( .A(ram[2971]), .B(n12850), .Y(n3228) );
  OAI21X1 U6180 ( .A(n12704), .B(n12850), .C(n3229), .Y(n7409) );
  NAND2X1 U6181 ( .A(ram[2972]), .B(n12850), .Y(n3229) );
  OAI21X1 U6182 ( .A(n12698), .B(n12850), .C(n3230), .Y(n7410) );
  NAND2X1 U6183 ( .A(ram[2973]), .B(n12850), .Y(n3230) );
  OAI21X1 U6184 ( .A(n12692), .B(n12850), .C(n3231), .Y(n7411) );
  NAND2X1 U6185 ( .A(ram[2974]), .B(n12850), .Y(n3231) );
  OAI21X1 U6186 ( .A(n12686), .B(n12850), .C(n3232), .Y(n7412) );
  NAND2X1 U6187 ( .A(ram[2975]), .B(n12850), .Y(n3232) );
  OAI21X1 U6189 ( .A(n12776), .B(n12849), .C(n3234), .Y(n7413) );
  NAND2X1 U6190 ( .A(ram[2976]), .B(n12849), .Y(n3234) );
  OAI21X1 U6191 ( .A(n12770), .B(n12849), .C(n3235), .Y(n7414) );
  NAND2X1 U6192 ( .A(ram[2977]), .B(n12849), .Y(n3235) );
  OAI21X1 U6193 ( .A(n12764), .B(n12849), .C(n3236), .Y(n7415) );
  NAND2X1 U6194 ( .A(ram[2978]), .B(n12849), .Y(n3236) );
  OAI21X1 U6195 ( .A(n12758), .B(n12849), .C(n3237), .Y(n7416) );
  NAND2X1 U6196 ( .A(ram[2979]), .B(n12849), .Y(n3237) );
  OAI21X1 U6197 ( .A(n12752), .B(n12849), .C(n3238), .Y(n7417) );
  NAND2X1 U6198 ( .A(ram[2980]), .B(n12849), .Y(n3238) );
  OAI21X1 U6199 ( .A(n12746), .B(n12849), .C(n3239), .Y(n7418) );
  NAND2X1 U6200 ( .A(ram[2981]), .B(n12849), .Y(n3239) );
  OAI21X1 U6201 ( .A(n12740), .B(n12849), .C(n3240), .Y(n7419) );
  NAND2X1 U6202 ( .A(ram[2982]), .B(n12849), .Y(n3240) );
  OAI21X1 U6203 ( .A(n12734), .B(n12849), .C(n3241), .Y(n7420) );
  NAND2X1 U6204 ( .A(ram[2983]), .B(n12849), .Y(n3241) );
  OAI21X1 U6205 ( .A(n12728), .B(n12849), .C(n3242), .Y(n7421) );
  NAND2X1 U6206 ( .A(ram[2984]), .B(n12849), .Y(n3242) );
  OAI21X1 U6207 ( .A(n12722), .B(n12849), .C(n3243), .Y(n7422) );
  NAND2X1 U6208 ( .A(ram[2985]), .B(n12849), .Y(n3243) );
  OAI21X1 U6209 ( .A(n12716), .B(n12849), .C(n3244), .Y(n7423) );
  NAND2X1 U6210 ( .A(ram[2986]), .B(n12849), .Y(n3244) );
  OAI21X1 U6211 ( .A(n12710), .B(n12849), .C(n3245), .Y(n7424) );
  NAND2X1 U6212 ( .A(ram[2987]), .B(n12849), .Y(n3245) );
  OAI21X1 U6213 ( .A(n12704), .B(n12849), .C(n3246), .Y(n7425) );
  NAND2X1 U6214 ( .A(ram[2988]), .B(n12849), .Y(n3246) );
  OAI21X1 U6215 ( .A(n12698), .B(n12849), .C(n3247), .Y(n7426) );
  NAND2X1 U6216 ( .A(ram[2989]), .B(n12849), .Y(n3247) );
  OAI21X1 U6217 ( .A(n12692), .B(n12849), .C(n3248), .Y(n7427) );
  NAND2X1 U6218 ( .A(ram[2990]), .B(n12849), .Y(n3248) );
  OAI21X1 U6219 ( .A(n12686), .B(n12849), .C(n3249), .Y(n7428) );
  NAND2X1 U6220 ( .A(ram[2991]), .B(n12849), .Y(n3249) );
  OAI21X1 U6222 ( .A(n12776), .B(n12848), .C(n3251), .Y(n7429) );
  NAND2X1 U6223 ( .A(ram[2992]), .B(n12848), .Y(n3251) );
  OAI21X1 U6224 ( .A(n12770), .B(n12848), .C(n3252), .Y(n7430) );
  NAND2X1 U6225 ( .A(ram[2993]), .B(n12848), .Y(n3252) );
  OAI21X1 U6226 ( .A(n12764), .B(n12848), .C(n3253), .Y(n7431) );
  NAND2X1 U6227 ( .A(ram[2994]), .B(n12848), .Y(n3253) );
  OAI21X1 U6228 ( .A(n12758), .B(n12848), .C(n3254), .Y(n7432) );
  NAND2X1 U6229 ( .A(ram[2995]), .B(n12848), .Y(n3254) );
  OAI21X1 U6230 ( .A(n12752), .B(n12848), .C(n3255), .Y(n7433) );
  NAND2X1 U6231 ( .A(ram[2996]), .B(n12848), .Y(n3255) );
  OAI21X1 U6232 ( .A(n12746), .B(n12848), .C(n3256), .Y(n7434) );
  NAND2X1 U6233 ( .A(ram[2997]), .B(n12848), .Y(n3256) );
  OAI21X1 U6234 ( .A(n12740), .B(n12848), .C(n3257), .Y(n7435) );
  NAND2X1 U6235 ( .A(ram[2998]), .B(n12848), .Y(n3257) );
  OAI21X1 U6236 ( .A(n12734), .B(n12848), .C(n3258), .Y(n7436) );
  NAND2X1 U6237 ( .A(ram[2999]), .B(n12848), .Y(n3258) );
  OAI21X1 U6238 ( .A(n12728), .B(n12848), .C(n3259), .Y(n7437) );
  NAND2X1 U6239 ( .A(ram[3000]), .B(n12848), .Y(n3259) );
  OAI21X1 U6240 ( .A(n12722), .B(n12848), .C(n3260), .Y(n7438) );
  NAND2X1 U6241 ( .A(ram[3001]), .B(n12848), .Y(n3260) );
  OAI21X1 U6242 ( .A(n12716), .B(n12848), .C(n3261), .Y(n7439) );
  NAND2X1 U6243 ( .A(ram[3002]), .B(n12848), .Y(n3261) );
  OAI21X1 U6244 ( .A(n12710), .B(n12848), .C(n3262), .Y(n7440) );
  NAND2X1 U6245 ( .A(ram[3003]), .B(n12848), .Y(n3262) );
  OAI21X1 U6246 ( .A(n12704), .B(n12848), .C(n3263), .Y(n7441) );
  NAND2X1 U6247 ( .A(ram[3004]), .B(n12848), .Y(n3263) );
  OAI21X1 U6248 ( .A(n12698), .B(n12848), .C(n3264), .Y(n7442) );
  NAND2X1 U6249 ( .A(ram[3005]), .B(n12848), .Y(n3264) );
  OAI21X1 U6250 ( .A(n12692), .B(n12848), .C(n3265), .Y(n7443) );
  NAND2X1 U6251 ( .A(ram[3006]), .B(n12848), .Y(n3265) );
  OAI21X1 U6252 ( .A(n12686), .B(n12848), .C(n3266), .Y(n7444) );
  NAND2X1 U6253 ( .A(ram[3007]), .B(n12848), .Y(n3266) );
  OAI21X1 U6255 ( .A(n12776), .B(n12847), .C(n3268), .Y(n7445) );
  NAND2X1 U6256 ( .A(ram[3008]), .B(n12847), .Y(n3268) );
  OAI21X1 U6257 ( .A(n12770), .B(n12847), .C(n3269), .Y(n7446) );
  NAND2X1 U6258 ( .A(ram[3009]), .B(n12847), .Y(n3269) );
  OAI21X1 U6259 ( .A(n12764), .B(n12847), .C(n3270), .Y(n7447) );
  NAND2X1 U6260 ( .A(ram[3010]), .B(n12847), .Y(n3270) );
  OAI21X1 U6261 ( .A(n12758), .B(n12847), .C(n3271), .Y(n7448) );
  NAND2X1 U6262 ( .A(ram[3011]), .B(n12847), .Y(n3271) );
  OAI21X1 U6263 ( .A(n12752), .B(n12847), .C(n3272), .Y(n7449) );
  NAND2X1 U6264 ( .A(ram[3012]), .B(n12847), .Y(n3272) );
  OAI21X1 U6265 ( .A(n12746), .B(n12847), .C(n3273), .Y(n7450) );
  NAND2X1 U6266 ( .A(ram[3013]), .B(n12847), .Y(n3273) );
  OAI21X1 U6267 ( .A(n12740), .B(n12847), .C(n3274), .Y(n7451) );
  NAND2X1 U6268 ( .A(ram[3014]), .B(n12847), .Y(n3274) );
  OAI21X1 U6269 ( .A(n12734), .B(n12847), .C(n3275), .Y(n7452) );
  NAND2X1 U6270 ( .A(ram[3015]), .B(n12847), .Y(n3275) );
  OAI21X1 U6271 ( .A(n12728), .B(n12847), .C(n3276), .Y(n7453) );
  NAND2X1 U6272 ( .A(ram[3016]), .B(n12847), .Y(n3276) );
  OAI21X1 U6273 ( .A(n12722), .B(n12847), .C(n3277), .Y(n7454) );
  NAND2X1 U6274 ( .A(ram[3017]), .B(n12847), .Y(n3277) );
  OAI21X1 U6275 ( .A(n12716), .B(n12847), .C(n3278), .Y(n7455) );
  NAND2X1 U6276 ( .A(ram[3018]), .B(n12847), .Y(n3278) );
  OAI21X1 U6277 ( .A(n12710), .B(n12847), .C(n3279), .Y(n7456) );
  NAND2X1 U6278 ( .A(ram[3019]), .B(n12847), .Y(n3279) );
  OAI21X1 U6279 ( .A(n12704), .B(n12847), .C(n3280), .Y(n7457) );
  NAND2X1 U6280 ( .A(ram[3020]), .B(n12847), .Y(n3280) );
  OAI21X1 U6281 ( .A(n12698), .B(n12847), .C(n3281), .Y(n7458) );
  NAND2X1 U6282 ( .A(ram[3021]), .B(n12847), .Y(n3281) );
  OAI21X1 U6283 ( .A(n12692), .B(n12847), .C(n3282), .Y(n7459) );
  NAND2X1 U6284 ( .A(ram[3022]), .B(n12847), .Y(n3282) );
  OAI21X1 U6285 ( .A(n12686), .B(n12847), .C(n3283), .Y(n7460) );
  NAND2X1 U6286 ( .A(ram[3023]), .B(n12847), .Y(n3283) );
  OAI21X1 U6288 ( .A(n12776), .B(n12846), .C(n3285), .Y(n7461) );
  NAND2X1 U6289 ( .A(ram[3024]), .B(n12846), .Y(n3285) );
  OAI21X1 U6290 ( .A(n12770), .B(n12846), .C(n3286), .Y(n7462) );
  NAND2X1 U6291 ( .A(ram[3025]), .B(n12846), .Y(n3286) );
  OAI21X1 U6292 ( .A(n12764), .B(n12846), .C(n3287), .Y(n7463) );
  NAND2X1 U6293 ( .A(ram[3026]), .B(n12846), .Y(n3287) );
  OAI21X1 U6294 ( .A(n12758), .B(n12846), .C(n3288), .Y(n7464) );
  NAND2X1 U6295 ( .A(ram[3027]), .B(n12846), .Y(n3288) );
  OAI21X1 U6296 ( .A(n12752), .B(n12846), .C(n3289), .Y(n7465) );
  NAND2X1 U6297 ( .A(ram[3028]), .B(n12846), .Y(n3289) );
  OAI21X1 U6298 ( .A(n12746), .B(n12846), .C(n3290), .Y(n7466) );
  NAND2X1 U6299 ( .A(ram[3029]), .B(n12846), .Y(n3290) );
  OAI21X1 U6300 ( .A(n12740), .B(n12846), .C(n3291), .Y(n7467) );
  NAND2X1 U6301 ( .A(ram[3030]), .B(n12846), .Y(n3291) );
  OAI21X1 U6302 ( .A(n12734), .B(n12846), .C(n3292), .Y(n7468) );
  NAND2X1 U6303 ( .A(ram[3031]), .B(n12846), .Y(n3292) );
  OAI21X1 U6304 ( .A(n12728), .B(n12846), .C(n3293), .Y(n7469) );
  NAND2X1 U6305 ( .A(ram[3032]), .B(n12846), .Y(n3293) );
  OAI21X1 U6306 ( .A(n12722), .B(n12846), .C(n3294), .Y(n7470) );
  NAND2X1 U6307 ( .A(ram[3033]), .B(n12846), .Y(n3294) );
  OAI21X1 U6308 ( .A(n12716), .B(n12846), .C(n3295), .Y(n7471) );
  NAND2X1 U6309 ( .A(ram[3034]), .B(n12846), .Y(n3295) );
  OAI21X1 U6310 ( .A(n12710), .B(n12846), .C(n3296), .Y(n7472) );
  NAND2X1 U6311 ( .A(ram[3035]), .B(n12846), .Y(n3296) );
  OAI21X1 U6312 ( .A(n12704), .B(n12846), .C(n3297), .Y(n7473) );
  NAND2X1 U6313 ( .A(ram[3036]), .B(n12846), .Y(n3297) );
  OAI21X1 U6314 ( .A(n12698), .B(n12846), .C(n3298), .Y(n7474) );
  NAND2X1 U6315 ( .A(ram[3037]), .B(n12846), .Y(n3298) );
  OAI21X1 U6316 ( .A(n12692), .B(n12846), .C(n3299), .Y(n7475) );
  NAND2X1 U6317 ( .A(ram[3038]), .B(n12846), .Y(n3299) );
  OAI21X1 U6318 ( .A(n12686), .B(n12846), .C(n3300), .Y(n7476) );
  NAND2X1 U6319 ( .A(ram[3039]), .B(n12846), .Y(n3300) );
  OAI21X1 U6321 ( .A(n12776), .B(n12845), .C(n3302), .Y(n7477) );
  NAND2X1 U6322 ( .A(ram[3040]), .B(n12845), .Y(n3302) );
  OAI21X1 U6323 ( .A(n12770), .B(n12845), .C(n3303), .Y(n7478) );
  NAND2X1 U6324 ( .A(ram[3041]), .B(n12845), .Y(n3303) );
  OAI21X1 U6325 ( .A(n12764), .B(n12845), .C(n3304), .Y(n7479) );
  NAND2X1 U6326 ( .A(ram[3042]), .B(n12845), .Y(n3304) );
  OAI21X1 U6327 ( .A(n12758), .B(n12845), .C(n3305), .Y(n7480) );
  NAND2X1 U6328 ( .A(ram[3043]), .B(n12845), .Y(n3305) );
  OAI21X1 U6329 ( .A(n12752), .B(n12845), .C(n3306), .Y(n7481) );
  NAND2X1 U6330 ( .A(ram[3044]), .B(n12845), .Y(n3306) );
  OAI21X1 U6331 ( .A(n12746), .B(n12845), .C(n3307), .Y(n7482) );
  NAND2X1 U6332 ( .A(ram[3045]), .B(n12845), .Y(n3307) );
  OAI21X1 U6333 ( .A(n12740), .B(n12845), .C(n3308), .Y(n7483) );
  NAND2X1 U6334 ( .A(ram[3046]), .B(n12845), .Y(n3308) );
  OAI21X1 U6335 ( .A(n12734), .B(n12845), .C(n3309), .Y(n7484) );
  NAND2X1 U6336 ( .A(ram[3047]), .B(n12845), .Y(n3309) );
  OAI21X1 U6337 ( .A(n12728), .B(n12845), .C(n3310), .Y(n7485) );
  NAND2X1 U6338 ( .A(ram[3048]), .B(n12845), .Y(n3310) );
  OAI21X1 U6339 ( .A(n12722), .B(n12845), .C(n3311), .Y(n7486) );
  NAND2X1 U6340 ( .A(ram[3049]), .B(n12845), .Y(n3311) );
  OAI21X1 U6341 ( .A(n12716), .B(n12845), .C(n3312), .Y(n7487) );
  NAND2X1 U6342 ( .A(ram[3050]), .B(n12845), .Y(n3312) );
  OAI21X1 U6343 ( .A(n12710), .B(n12845), .C(n3313), .Y(n7488) );
  NAND2X1 U6344 ( .A(ram[3051]), .B(n12845), .Y(n3313) );
  OAI21X1 U6345 ( .A(n12704), .B(n12845), .C(n3314), .Y(n7489) );
  NAND2X1 U6346 ( .A(ram[3052]), .B(n12845), .Y(n3314) );
  OAI21X1 U6347 ( .A(n12698), .B(n12845), .C(n3315), .Y(n7490) );
  NAND2X1 U6348 ( .A(ram[3053]), .B(n12845), .Y(n3315) );
  OAI21X1 U6349 ( .A(n12692), .B(n12845), .C(n3316), .Y(n7491) );
  NAND2X1 U6350 ( .A(ram[3054]), .B(n12845), .Y(n3316) );
  OAI21X1 U6351 ( .A(n12686), .B(n12845), .C(n3317), .Y(n7492) );
  NAND2X1 U6352 ( .A(ram[3055]), .B(n12845), .Y(n3317) );
  OAI21X1 U6354 ( .A(n12776), .B(n12844), .C(n3319), .Y(n7493) );
  NAND2X1 U6355 ( .A(ram[3056]), .B(n12844), .Y(n3319) );
  OAI21X1 U6356 ( .A(n12770), .B(n12844), .C(n3320), .Y(n7494) );
  NAND2X1 U6357 ( .A(ram[3057]), .B(n12844), .Y(n3320) );
  OAI21X1 U6358 ( .A(n12764), .B(n12844), .C(n3321), .Y(n7495) );
  NAND2X1 U6359 ( .A(ram[3058]), .B(n12844), .Y(n3321) );
  OAI21X1 U6360 ( .A(n12758), .B(n12844), .C(n3322), .Y(n7496) );
  NAND2X1 U6361 ( .A(ram[3059]), .B(n12844), .Y(n3322) );
  OAI21X1 U6362 ( .A(n12752), .B(n12844), .C(n3323), .Y(n7497) );
  NAND2X1 U6363 ( .A(ram[3060]), .B(n12844), .Y(n3323) );
  OAI21X1 U6364 ( .A(n12746), .B(n12844), .C(n3324), .Y(n7498) );
  NAND2X1 U6365 ( .A(ram[3061]), .B(n12844), .Y(n3324) );
  OAI21X1 U6366 ( .A(n12740), .B(n12844), .C(n3325), .Y(n7499) );
  NAND2X1 U6367 ( .A(ram[3062]), .B(n12844), .Y(n3325) );
  OAI21X1 U6368 ( .A(n12734), .B(n12844), .C(n3326), .Y(n7500) );
  NAND2X1 U6369 ( .A(ram[3063]), .B(n12844), .Y(n3326) );
  OAI21X1 U6370 ( .A(n12728), .B(n12844), .C(n3327), .Y(n7501) );
  NAND2X1 U6371 ( .A(ram[3064]), .B(n12844), .Y(n3327) );
  OAI21X1 U6372 ( .A(n12722), .B(n12844), .C(n3328), .Y(n7502) );
  NAND2X1 U6373 ( .A(ram[3065]), .B(n12844), .Y(n3328) );
  OAI21X1 U6374 ( .A(n12716), .B(n12844), .C(n3329), .Y(n7503) );
  NAND2X1 U6375 ( .A(ram[3066]), .B(n12844), .Y(n3329) );
  OAI21X1 U6376 ( .A(n12710), .B(n12844), .C(n3330), .Y(n7504) );
  NAND2X1 U6377 ( .A(ram[3067]), .B(n12844), .Y(n3330) );
  OAI21X1 U6378 ( .A(n12704), .B(n12844), .C(n3331), .Y(n7505) );
  NAND2X1 U6379 ( .A(ram[3068]), .B(n12844), .Y(n3331) );
  OAI21X1 U6380 ( .A(n12698), .B(n12844), .C(n3332), .Y(n7506) );
  NAND2X1 U6381 ( .A(ram[3069]), .B(n12844), .Y(n3332) );
  OAI21X1 U6382 ( .A(n12692), .B(n12844), .C(n3333), .Y(n7507) );
  NAND2X1 U6383 ( .A(ram[3070]), .B(n12844), .Y(n3333) );
  OAI21X1 U6384 ( .A(n12686), .B(n12844), .C(n3334), .Y(n7508) );
  NAND2X1 U6385 ( .A(ram[3071]), .B(n12844), .Y(n3334) );
  NAND3X1 U6387 ( .A(n1149), .B(mem_write_en), .C(n2516), .Y(n3335) );
  AND2X1 U6388 ( .A(mem_access_addr[7]), .B(n13039), .Y(n2516) );
  OAI21X1 U6389 ( .A(n12776), .B(n12843), .C(n3337), .Y(n7509) );
  NAND2X1 U6390 ( .A(ram[3072]), .B(n12843), .Y(n3337) );
  OAI21X1 U6391 ( .A(n12770), .B(n12843), .C(n3338), .Y(n7510) );
  NAND2X1 U6392 ( .A(ram[3073]), .B(n12843), .Y(n3338) );
  OAI21X1 U6393 ( .A(n12764), .B(n12843), .C(n3339), .Y(n7511) );
  NAND2X1 U6394 ( .A(ram[3074]), .B(n12843), .Y(n3339) );
  OAI21X1 U6395 ( .A(n12758), .B(n12843), .C(n3340), .Y(n7512) );
  NAND2X1 U6396 ( .A(ram[3075]), .B(n12843), .Y(n3340) );
  OAI21X1 U6397 ( .A(n12752), .B(n12843), .C(n3341), .Y(n7513) );
  NAND2X1 U6398 ( .A(ram[3076]), .B(n12843), .Y(n3341) );
  OAI21X1 U6399 ( .A(n12746), .B(n12843), .C(n3342), .Y(n7514) );
  NAND2X1 U6400 ( .A(ram[3077]), .B(n12843), .Y(n3342) );
  OAI21X1 U6401 ( .A(n12740), .B(n12843), .C(n3343), .Y(n7515) );
  NAND2X1 U6402 ( .A(ram[3078]), .B(n12843), .Y(n3343) );
  OAI21X1 U6403 ( .A(n12734), .B(n12843), .C(n3344), .Y(n7516) );
  NAND2X1 U6404 ( .A(ram[3079]), .B(n12843), .Y(n3344) );
  OAI21X1 U6405 ( .A(n12728), .B(n12843), .C(n3345), .Y(n7517) );
  NAND2X1 U6406 ( .A(ram[3080]), .B(n12843), .Y(n3345) );
  OAI21X1 U6407 ( .A(n12722), .B(n12843), .C(n3346), .Y(n7518) );
  NAND2X1 U6408 ( .A(ram[3081]), .B(n12843), .Y(n3346) );
  OAI21X1 U6409 ( .A(n12716), .B(n12843), .C(n3347), .Y(n7519) );
  NAND2X1 U6410 ( .A(ram[3082]), .B(n12843), .Y(n3347) );
  OAI21X1 U6411 ( .A(n12710), .B(n12843), .C(n3348), .Y(n7520) );
  NAND2X1 U6412 ( .A(ram[3083]), .B(n12843), .Y(n3348) );
  OAI21X1 U6413 ( .A(n12704), .B(n12843), .C(n3349), .Y(n7521) );
  NAND2X1 U6414 ( .A(ram[3084]), .B(n12843), .Y(n3349) );
  OAI21X1 U6415 ( .A(n12698), .B(n12843), .C(n3350), .Y(n7522) );
  NAND2X1 U6416 ( .A(ram[3085]), .B(n12843), .Y(n3350) );
  OAI21X1 U6417 ( .A(n12692), .B(n12843), .C(n3351), .Y(n7523) );
  NAND2X1 U6418 ( .A(ram[3086]), .B(n12843), .Y(n3351) );
  OAI21X1 U6419 ( .A(n12686), .B(n12843), .C(n3352), .Y(n7524) );
  NAND2X1 U6420 ( .A(ram[3087]), .B(n12843), .Y(n3352) );
  OAI21X1 U6422 ( .A(n12776), .B(n12842), .C(n3354), .Y(n7525) );
  NAND2X1 U6423 ( .A(ram[3088]), .B(n12842), .Y(n3354) );
  OAI21X1 U6424 ( .A(n12770), .B(n12842), .C(n3355), .Y(n7526) );
  NAND2X1 U6425 ( .A(ram[3089]), .B(n12842), .Y(n3355) );
  OAI21X1 U6426 ( .A(n12764), .B(n12842), .C(n3356), .Y(n7527) );
  NAND2X1 U6427 ( .A(ram[3090]), .B(n12842), .Y(n3356) );
  OAI21X1 U6428 ( .A(n12758), .B(n12842), .C(n3357), .Y(n7528) );
  NAND2X1 U6429 ( .A(ram[3091]), .B(n12842), .Y(n3357) );
  OAI21X1 U6430 ( .A(n12752), .B(n12842), .C(n3358), .Y(n7529) );
  NAND2X1 U6431 ( .A(ram[3092]), .B(n12842), .Y(n3358) );
  OAI21X1 U6432 ( .A(n12746), .B(n12842), .C(n3359), .Y(n7530) );
  NAND2X1 U6433 ( .A(ram[3093]), .B(n12842), .Y(n3359) );
  OAI21X1 U6434 ( .A(n12740), .B(n12842), .C(n3360), .Y(n7531) );
  NAND2X1 U6435 ( .A(ram[3094]), .B(n12842), .Y(n3360) );
  OAI21X1 U6436 ( .A(n12734), .B(n12842), .C(n3361), .Y(n7532) );
  NAND2X1 U6437 ( .A(ram[3095]), .B(n12842), .Y(n3361) );
  OAI21X1 U6438 ( .A(n12728), .B(n12842), .C(n3362), .Y(n7533) );
  NAND2X1 U6439 ( .A(ram[3096]), .B(n12842), .Y(n3362) );
  OAI21X1 U6440 ( .A(n12722), .B(n12842), .C(n3363), .Y(n7534) );
  NAND2X1 U6441 ( .A(ram[3097]), .B(n12842), .Y(n3363) );
  OAI21X1 U6442 ( .A(n12716), .B(n12842), .C(n3364), .Y(n7535) );
  NAND2X1 U6443 ( .A(ram[3098]), .B(n12842), .Y(n3364) );
  OAI21X1 U6444 ( .A(n12710), .B(n12842), .C(n3365), .Y(n7536) );
  NAND2X1 U6445 ( .A(ram[3099]), .B(n12842), .Y(n3365) );
  OAI21X1 U6446 ( .A(n12704), .B(n12842), .C(n3366), .Y(n7537) );
  NAND2X1 U6447 ( .A(ram[3100]), .B(n12842), .Y(n3366) );
  OAI21X1 U6448 ( .A(n12698), .B(n12842), .C(n3367), .Y(n7538) );
  NAND2X1 U6449 ( .A(ram[3101]), .B(n12842), .Y(n3367) );
  OAI21X1 U6450 ( .A(n12692), .B(n12842), .C(n3368), .Y(n7539) );
  NAND2X1 U6451 ( .A(ram[3102]), .B(n12842), .Y(n3368) );
  OAI21X1 U6452 ( .A(n12686), .B(n12842), .C(n3369), .Y(n7540) );
  NAND2X1 U6453 ( .A(ram[3103]), .B(n12842), .Y(n3369) );
  OAI21X1 U6455 ( .A(n12776), .B(n12841), .C(n3371), .Y(n7541) );
  NAND2X1 U6456 ( .A(ram[3104]), .B(n12841), .Y(n3371) );
  OAI21X1 U6457 ( .A(n12770), .B(n12841), .C(n3372), .Y(n7542) );
  NAND2X1 U6458 ( .A(ram[3105]), .B(n12841), .Y(n3372) );
  OAI21X1 U6459 ( .A(n12764), .B(n12841), .C(n3373), .Y(n7543) );
  NAND2X1 U6460 ( .A(ram[3106]), .B(n12841), .Y(n3373) );
  OAI21X1 U6461 ( .A(n12758), .B(n12841), .C(n3374), .Y(n7544) );
  NAND2X1 U6462 ( .A(ram[3107]), .B(n12841), .Y(n3374) );
  OAI21X1 U6463 ( .A(n12752), .B(n12841), .C(n3375), .Y(n7545) );
  NAND2X1 U6464 ( .A(ram[3108]), .B(n12841), .Y(n3375) );
  OAI21X1 U6465 ( .A(n12746), .B(n12841), .C(n3376), .Y(n7546) );
  NAND2X1 U6466 ( .A(ram[3109]), .B(n12841), .Y(n3376) );
  OAI21X1 U6467 ( .A(n12740), .B(n12841), .C(n3377), .Y(n7547) );
  NAND2X1 U6468 ( .A(ram[3110]), .B(n12841), .Y(n3377) );
  OAI21X1 U6469 ( .A(n12734), .B(n12841), .C(n3378), .Y(n7548) );
  NAND2X1 U6470 ( .A(ram[3111]), .B(n12841), .Y(n3378) );
  OAI21X1 U6471 ( .A(n12728), .B(n12841), .C(n3379), .Y(n7549) );
  NAND2X1 U6472 ( .A(ram[3112]), .B(n12841), .Y(n3379) );
  OAI21X1 U6473 ( .A(n12722), .B(n12841), .C(n3380), .Y(n7550) );
  NAND2X1 U6474 ( .A(ram[3113]), .B(n12841), .Y(n3380) );
  OAI21X1 U6475 ( .A(n12716), .B(n12841), .C(n3381), .Y(n7551) );
  NAND2X1 U6476 ( .A(ram[3114]), .B(n12841), .Y(n3381) );
  OAI21X1 U6477 ( .A(n12710), .B(n12841), .C(n3382), .Y(n7552) );
  NAND2X1 U6478 ( .A(ram[3115]), .B(n12841), .Y(n3382) );
  OAI21X1 U6479 ( .A(n12704), .B(n12841), .C(n3383), .Y(n7553) );
  NAND2X1 U6480 ( .A(ram[3116]), .B(n12841), .Y(n3383) );
  OAI21X1 U6481 ( .A(n12698), .B(n12841), .C(n3384), .Y(n7554) );
  NAND2X1 U6482 ( .A(ram[3117]), .B(n12841), .Y(n3384) );
  OAI21X1 U6483 ( .A(n12692), .B(n12841), .C(n3385), .Y(n7555) );
  NAND2X1 U6484 ( .A(ram[3118]), .B(n12841), .Y(n3385) );
  OAI21X1 U6485 ( .A(n12686), .B(n12841), .C(n3386), .Y(n7556) );
  NAND2X1 U6486 ( .A(ram[3119]), .B(n12841), .Y(n3386) );
  OAI21X1 U6488 ( .A(n12777), .B(n12840), .C(n3388), .Y(n7557) );
  NAND2X1 U6489 ( .A(ram[3120]), .B(n12840), .Y(n3388) );
  OAI21X1 U6490 ( .A(n12771), .B(n12840), .C(n3389), .Y(n7558) );
  NAND2X1 U6491 ( .A(ram[3121]), .B(n12840), .Y(n3389) );
  OAI21X1 U6492 ( .A(n12765), .B(n12840), .C(n3390), .Y(n7559) );
  NAND2X1 U6493 ( .A(ram[3122]), .B(n12840), .Y(n3390) );
  OAI21X1 U6494 ( .A(n12759), .B(n12840), .C(n3391), .Y(n7560) );
  NAND2X1 U6495 ( .A(ram[3123]), .B(n12840), .Y(n3391) );
  OAI21X1 U6496 ( .A(n12753), .B(n12840), .C(n3392), .Y(n7561) );
  NAND2X1 U6497 ( .A(ram[3124]), .B(n12840), .Y(n3392) );
  OAI21X1 U6498 ( .A(n12747), .B(n12840), .C(n3393), .Y(n7562) );
  NAND2X1 U6499 ( .A(ram[3125]), .B(n12840), .Y(n3393) );
  OAI21X1 U6500 ( .A(n12741), .B(n12840), .C(n3394), .Y(n7563) );
  NAND2X1 U6501 ( .A(ram[3126]), .B(n12840), .Y(n3394) );
  OAI21X1 U6502 ( .A(n12735), .B(n12840), .C(n3395), .Y(n7564) );
  NAND2X1 U6503 ( .A(ram[3127]), .B(n12840), .Y(n3395) );
  OAI21X1 U6504 ( .A(n12729), .B(n12840), .C(n3396), .Y(n7565) );
  NAND2X1 U6505 ( .A(ram[3128]), .B(n12840), .Y(n3396) );
  OAI21X1 U6506 ( .A(n12723), .B(n12840), .C(n3397), .Y(n7566) );
  NAND2X1 U6507 ( .A(ram[3129]), .B(n12840), .Y(n3397) );
  OAI21X1 U6508 ( .A(n12717), .B(n12840), .C(n3398), .Y(n7567) );
  NAND2X1 U6509 ( .A(ram[3130]), .B(n12840), .Y(n3398) );
  OAI21X1 U6510 ( .A(n12711), .B(n12840), .C(n3399), .Y(n7568) );
  NAND2X1 U6511 ( .A(ram[3131]), .B(n12840), .Y(n3399) );
  OAI21X1 U6512 ( .A(n12705), .B(n12840), .C(n3400), .Y(n7569) );
  NAND2X1 U6513 ( .A(ram[3132]), .B(n12840), .Y(n3400) );
  OAI21X1 U6514 ( .A(n12699), .B(n12840), .C(n3401), .Y(n7570) );
  NAND2X1 U6515 ( .A(ram[3133]), .B(n12840), .Y(n3401) );
  OAI21X1 U6516 ( .A(n12693), .B(n12840), .C(n3402), .Y(n7571) );
  NAND2X1 U6517 ( .A(ram[3134]), .B(n12840), .Y(n3402) );
  OAI21X1 U6518 ( .A(n12687), .B(n12840), .C(n3403), .Y(n7572) );
  NAND2X1 U6519 ( .A(ram[3135]), .B(n12840), .Y(n3403) );
  OAI21X1 U6521 ( .A(n12777), .B(n12839), .C(n3405), .Y(n7573) );
  NAND2X1 U6522 ( .A(ram[3136]), .B(n12839), .Y(n3405) );
  OAI21X1 U6523 ( .A(n12771), .B(n12839), .C(n3406), .Y(n7574) );
  NAND2X1 U6524 ( .A(ram[3137]), .B(n12839), .Y(n3406) );
  OAI21X1 U6525 ( .A(n12765), .B(n12839), .C(n3407), .Y(n7575) );
  NAND2X1 U6526 ( .A(ram[3138]), .B(n12839), .Y(n3407) );
  OAI21X1 U6527 ( .A(n12759), .B(n12839), .C(n3408), .Y(n7576) );
  NAND2X1 U6528 ( .A(ram[3139]), .B(n12839), .Y(n3408) );
  OAI21X1 U6529 ( .A(n12753), .B(n12839), .C(n3409), .Y(n7577) );
  NAND2X1 U6530 ( .A(ram[3140]), .B(n12839), .Y(n3409) );
  OAI21X1 U6531 ( .A(n12747), .B(n12839), .C(n3410), .Y(n7578) );
  NAND2X1 U6532 ( .A(ram[3141]), .B(n12839), .Y(n3410) );
  OAI21X1 U6533 ( .A(n12741), .B(n12839), .C(n3411), .Y(n7579) );
  NAND2X1 U6534 ( .A(ram[3142]), .B(n12839), .Y(n3411) );
  OAI21X1 U6535 ( .A(n12735), .B(n12839), .C(n3412), .Y(n7580) );
  NAND2X1 U6536 ( .A(ram[3143]), .B(n12839), .Y(n3412) );
  OAI21X1 U6537 ( .A(n12729), .B(n12839), .C(n3413), .Y(n7581) );
  NAND2X1 U6538 ( .A(ram[3144]), .B(n12839), .Y(n3413) );
  OAI21X1 U6539 ( .A(n12723), .B(n12839), .C(n3414), .Y(n7582) );
  NAND2X1 U6540 ( .A(ram[3145]), .B(n12839), .Y(n3414) );
  OAI21X1 U6541 ( .A(n12717), .B(n12839), .C(n3415), .Y(n7583) );
  NAND2X1 U6542 ( .A(ram[3146]), .B(n12839), .Y(n3415) );
  OAI21X1 U6543 ( .A(n12711), .B(n12839), .C(n3416), .Y(n7584) );
  NAND2X1 U6544 ( .A(ram[3147]), .B(n12839), .Y(n3416) );
  OAI21X1 U6545 ( .A(n12705), .B(n12839), .C(n3417), .Y(n7585) );
  NAND2X1 U6546 ( .A(ram[3148]), .B(n12839), .Y(n3417) );
  OAI21X1 U6547 ( .A(n12699), .B(n12839), .C(n3418), .Y(n7586) );
  NAND2X1 U6548 ( .A(ram[3149]), .B(n12839), .Y(n3418) );
  OAI21X1 U6549 ( .A(n12693), .B(n12839), .C(n3419), .Y(n7587) );
  NAND2X1 U6550 ( .A(ram[3150]), .B(n12839), .Y(n3419) );
  OAI21X1 U6551 ( .A(n12687), .B(n12839), .C(n3420), .Y(n7588) );
  NAND2X1 U6552 ( .A(ram[3151]), .B(n12839), .Y(n3420) );
  OAI21X1 U6554 ( .A(n12777), .B(n12838), .C(n3422), .Y(n7589) );
  NAND2X1 U6555 ( .A(ram[3152]), .B(n12838), .Y(n3422) );
  OAI21X1 U6556 ( .A(n12771), .B(n12838), .C(n3423), .Y(n7590) );
  NAND2X1 U6557 ( .A(ram[3153]), .B(n12838), .Y(n3423) );
  OAI21X1 U6558 ( .A(n12765), .B(n12838), .C(n3424), .Y(n7591) );
  NAND2X1 U6559 ( .A(ram[3154]), .B(n12838), .Y(n3424) );
  OAI21X1 U6560 ( .A(n12759), .B(n12838), .C(n3425), .Y(n7592) );
  NAND2X1 U6561 ( .A(ram[3155]), .B(n12838), .Y(n3425) );
  OAI21X1 U6562 ( .A(n12753), .B(n12838), .C(n3426), .Y(n7593) );
  NAND2X1 U6563 ( .A(ram[3156]), .B(n12838), .Y(n3426) );
  OAI21X1 U6564 ( .A(n12747), .B(n12838), .C(n3427), .Y(n7594) );
  NAND2X1 U6565 ( .A(ram[3157]), .B(n12838), .Y(n3427) );
  OAI21X1 U6566 ( .A(n12741), .B(n12838), .C(n3428), .Y(n7595) );
  NAND2X1 U6567 ( .A(ram[3158]), .B(n12838), .Y(n3428) );
  OAI21X1 U6568 ( .A(n12735), .B(n12838), .C(n3429), .Y(n7596) );
  NAND2X1 U6569 ( .A(ram[3159]), .B(n12838), .Y(n3429) );
  OAI21X1 U6570 ( .A(n12729), .B(n12838), .C(n3430), .Y(n7597) );
  NAND2X1 U6571 ( .A(ram[3160]), .B(n12838), .Y(n3430) );
  OAI21X1 U6572 ( .A(n12723), .B(n12838), .C(n3431), .Y(n7598) );
  NAND2X1 U6573 ( .A(ram[3161]), .B(n12838), .Y(n3431) );
  OAI21X1 U6574 ( .A(n12717), .B(n12838), .C(n3432), .Y(n7599) );
  NAND2X1 U6575 ( .A(ram[3162]), .B(n12838), .Y(n3432) );
  OAI21X1 U6576 ( .A(n12711), .B(n12838), .C(n3433), .Y(n7600) );
  NAND2X1 U6577 ( .A(ram[3163]), .B(n12838), .Y(n3433) );
  OAI21X1 U6578 ( .A(n12705), .B(n12838), .C(n3434), .Y(n7601) );
  NAND2X1 U6579 ( .A(ram[3164]), .B(n12838), .Y(n3434) );
  OAI21X1 U6580 ( .A(n12699), .B(n12838), .C(n3435), .Y(n7602) );
  NAND2X1 U6581 ( .A(ram[3165]), .B(n12838), .Y(n3435) );
  OAI21X1 U6582 ( .A(n12693), .B(n12838), .C(n3436), .Y(n7603) );
  NAND2X1 U6583 ( .A(ram[3166]), .B(n12838), .Y(n3436) );
  OAI21X1 U6584 ( .A(n12687), .B(n12838), .C(n3437), .Y(n7604) );
  NAND2X1 U6585 ( .A(ram[3167]), .B(n12838), .Y(n3437) );
  OAI21X1 U6587 ( .A(n12777), .B(n12837), .C(n3439), .Y(n7605) );
  NAND2X1 U6588 ( .A(ram[3168]), .B(n12837), .Y(n3439) );
  OAI21X1 U6589 ( .A(n12771), .B(n12837), .C(n3440), .Y(n7606) );
  NAND2X1 U6590 ( .A(ram[3169]), .B(n12837), .Y(n3440) );
  OAI21X1 U6591 ( .A(n12765), .B(n12837), .C(n3441), .Y(n7607) );
  NAND2X1 U6592 ( .A(ram[3170]), .B(n12837), .Y(n3441) );
  OAI21X1 U6593 ( .A(n12759), .B(n12837), .C(n3442), .Y(n7608) );
  NAND2X1 U6594 ( .A(ram[3171]), .B(n12837), .Y(n3442) );
  OAI21X1 U6595 ( .A(n12753), .B(n12837), .C(n3443), .Y(n7609) );
  NAND2X1 U6596 ( .A(ram[3172]), .B(n12837), .Y(n3443) );
  OAI21X1 U6597 ( .A(n12747), .B(n12837), .C(n3444), .Y(n7610) );
  NAND2X1 U6598 ( .A(ram[3173]), .B(n12837), .Y(n3444) );
  OAI21X1 U6599 ( .A(n12741), .B(n12837), .C(n3445), .Y(n7611) );
  NAND2X1 U6600 ( .A(ram[3174]), .B(n12837), .Y(n3445) );
  OAI21X1 U6601 ( .A(n12735), .B(n12837), .C(n3446), .Y(n7612) );
  NAND2X1 U6602 ( .A(ram[3175]), .B(n12837), .Y(n3446) );
  OAI21X1 U6603 ( .A(n12729), .B(n12837), .C(n3447), .Y(n7613) );
  NAND2X1 U6604 ( .A(ram[3176]), .B(n12837), .Y(n3447) );
  OAI21X1 U6605 ( .A(n12723), .B(n12837), .C(n3448), .Y(n7614) );
  NAND2X1 U6606 ( .A(ram[3177]), .B(n12837), .Y(n3448) );
  OAI21X1 U6607 ( .A(n12717), .B(n12837), .C(n3449), .Y(n7615) );
  NAND2X1 U6608 ( .A(ram[3178]), .B(n12837), .Y(n3449) );
  OAI21X1 U6609 ( .A(n12711), .B(n12837), .C(n3450), .Y(n7616) );
  NAND2X1 U6610 ( .A(ram[3179]), .B(n12837), .Y(n3450) );
  OAI21X1 U6611 ( .A(n12705), .B(n12837), .C(n3451), .Y(n7617) );
  NAND2X1 U6612 ( .A(ram[3180]), .B(n12837), .Y(n3451) );
  OAI21X1 U6613 ( .A(n12699), .B(n12837), .C(n3452), .Y(n7618) );
  NAND2X1 U6614 ( .A(ram[3181]), .B(n12837), .Y(n3452) );
  OAI21X1 U6615 ( .A(n12693), .B(n12837), .C(n3453), .Y(n7619) );
  NAND2X1 U6616 ( .A(ram[3182]), .B(n12837), .Y(n3453) );
  OAI21X1 U6617 ( .A(n12687), .B(n12837), .C(n3454), .Y(n7620) );
  NAND2X1 U6618 ( .A(ram[3183]), .B(n12837), .Y(n3454) );
  OAI21X1 U6620 ( .A(n12777), .B(n12836), .C(n3456), .Y(n7621) );
  NAND2X1 U6621 ( .A(ram[3184]), .B(n12836), .Y(n3456) );
  OAI21X1 U6622 ( .A(n12771), .B(n12836), .C(n3457), .Y(n7622) );
  NAND2X1 U6623 ( .A(ram[3185]), .B(n12836), .Y(n3457) );
  OAI21X1 U6624 ( .A(n12765), .B(n12836), .C(n3458), .Y(n7623) );
  NAND2X1 U6625 ( .A(ram[3186]), .B(n12836), .Y(n3458) );
  OAI21X1 U6626 ( .A(n12759), .B(n12836), .C(n3459), .Y(n7624) );
  NAND2X1 U6627 ( .A(ram[3187]), .B(n12836), .Y(n3459) );
  OAI21X1 U6628 ( .A(n12753), .B(n12836), .C(n3460), .Y(n7625) );
  NAND2X1 U6629 ( .A(ram[3188]), .B(n12836), .Y(n3460) );
  OAI21X1 U6630 ( .A(n12747), .B(n12836), .C(n3461), .Y(n7626) );
  NAND2X1 U6631 ( .A(ram[3189]), .B(n12836), .Y(n3461) );
  OAI21X1 U6632 ( .A(n12741), .B(n12836), .C(n3462), .Y(n7627) );
  NAND2X1 U6633 ( .A(ram[3190]), .B(n12836), .Y(n3462) );
  OAI21X1 U6634 ( .A(n12735), .B(n12836), .C(n3463), .Y(n7628) );
  NAND2X1 U6635 ( .A(ram[3191]), .B(n12836), .Y(n3463) );
  OAI21X1 U6636 ( .A(n12729), .B(n12836), .C(n3464), .Y(n7629) );
  NAND2X1 U6637 ( .A(ram[3192]), .B(n12836), .Y(n3464) );
  OAI21X1 U6638 ( .A(n12723), .B(n12836), .C(n3465), .Y(n7630) );
  NAND2X1 U6639 ( .A(ram[3193]), .B(n12836), .Y(n3465) );
  OAI21X1 U6640 ( .A(n12717), .B(n12836), .C(n3466), .Y(n7631) );
  NAND2X1 U6641 ( .A(ram[3194]), .B(n12836), .Y(n3466) );
  OAI21X1 U6642 ( .A(n12711), .B(n12836), .C(n3467), .Y(n7632) );
  NAND2X1 U6643 ( .A(ram[3195]), .B(n12836), .Y(n3467) );
  OAI21X1 U6644 ( .A(n12705), .B(n12836), .C(n3468), .Y(n7633) );
  NAND2X1 U6645 ( .A(ram[3196]), .B(n12836), .Y(n3468) );
  OAI21X1 U6646 ( .A(n12699), .B(n12836), .C(n3469), .Y(n7634) );
  NAND2X1 U6647 ( .A(ram[3197]), .B(n12836), .Y(n3469) );
  OAI21X1 U6648 ( .A(n12693), .B(n12836), .C(n3470), .Y(n7635) );
  NAND2X1 U6649 ( .A(ram[3198]), .B(n12836), .Y(n3470) );
  OAI21X1 U6650 ( .A(n12687), .B(n12836), .C(n3471), .Y(n7636) );
  NAND2X1 U6651 ( .A(ram[3199]), .B(n12836), .Y(n3471) );
  OAI21X1 U6653 ( .A(n12777), .B(n12835), .C(n3473), .Y(n7637) );
  NAND2X1 U6654 ( .A(ram[3200]), .B(n12835), .Y(n3473) );
  OAI21X1 U6655 ( .A(n12771), .B(n12835), .C(n3474), .Y(n7638) );
  NAND2X1 U6656 ( .A(ram[3201]), .B(n12835), .Y(n3474) );
  OAI21X1 U6657 ( .A(n12765), .B(n12835), .C(n3475), .Y(n7639) );
  NAND2X1 U6658 ( .A(ram[3202]), .B(n12835), .Y(n3475) );
  OAI21X1 U6659 ( .A(n12759), .B(n12835), .C(n3476), .Y(n7640) );
  NAND2X1 U6660 ( .A(ram[3203]), .B(n12835), .Y(n3476) );
  OAI21X1 U6661 ( .A(n12753), .B(n12835), .C(n3477), .Y(n7641) );
  NAND2X1 U6662 ( .A(ram[3204]), .B(n12835), .Y(n3477) );
  OAI21X1 U6663 ( .A(n12747), .B(n12835), .C(n3478), .Y(n7642) );
  NAND2X1 U6664 ( .A(ram[3205]), .B(n12835), .Y(n3478) );
  OAI21X1 U6665 ( .A(n12741), .B(n12835), .C(n3479), .Y(n7643) );
  NAND2X1 U6666 ( .A(ram[3206]), .B(n12835), .Y(n3479) );
  OAI21X1 U6667 ( .A(n12735), .B(n12835), .C(n3480), .Y(n7644) );
  NAND2X1 U6668 ( .A(ram[3207]), .B(n12835), .Y(n3480) );
  OAI21X1 U6669 ( .A(n12729), .B(n12835), .C(n3481), .Y(n7645) );
  NAND2X1 U6670 ( .A(ram[3208]), .B(n12835), .Y(n3481) );
  OAI21X1 U6671 ( .A(n12723), .B(n12835), .C(n3482), .Y(n7646) );
  NAND2X1 U6672 ( .A(ram[3209]), .B(n12835), .Y(n3482) );
  OAI21X1 U6673 ( .A(n12717), .B(n12835), .C(n3483), .Y(n7647) );
  NAND2X1 U6674 ( .A(ram[3210]), .B(n12835), .Y(n3483) );
  OAI21X1 U6675 ( .A(n12711), .B(n12835), .C(n3484), .Y(n7648) );
  NAND2X1 U6676 ( .A(ram[3211]), .B(n12835), .Y(n3484) );
  OAI21X1 U6677 ( .A(n12705), .B(n12835), .C(n3485), .Y(n7649) );
  NAND2X1 U6678 ( .A(ram[3212]), .B(n12835), .Y(n3485) );
  OAI21X1 U6679 ( .A(n12699), .B(n12835), .C(n3486), .Y(n7650) );
  NAND2X1 U6680 ( .A(ram[3213]), .B(n12835), .Y(n3486) );
  OAI21X1 U6681 ( .A(n12693), .B(n12835), .C(n3487), .Y(n7651) );
  NAND2X1 U6682 ( .A(ram[3214]), .B(n12835), .Y(n3487) );
  OAI21X1 U6683 ( .A(n12687), .B(n12835), .C(n3488), .Y(n7652) );
  NAND2X1 U6684 ( .A(ram[3215]), .B(n12835), .Y(n3488) );
  OAI21X1 U6686 ( .A(n12777), .B(n12834), .C(n3490), .Y(n7653) );
  NAND2X1 U6687 ( .A(ram[3216]), .B(n12834), .Y(n3490) );
  OAI21X1 U6688 ( .A(n12771), .B(n12834), .C(n3491), .Y(n7654) );
  NAND2X1 U6689 ( .A(ram[3217]), .B(n12834), .Y(n3491) );
  OAI21X1 U6690 ( .A(n12765), .B(n12834), .C(n3492), .Y(n7655) );
  NAND2X1 U6691 ( .A(ram[3218]), .B(n12834), .Y(n3492) );
  OAI21X1 U6692 ( .A(n12759), .B(n12834), .C(n3493), .Y(n7656) );
  NAND2X1 U6693 ( .A(ram[3219]), .B(n12834), .Y(n3493) );
  OAI21X1 U6694 ( .A(n12753), .B(n12834), .C(n3494), .Y(n7657) );
  NAND2X1 U6695 ( .A(ram[3220]), .B(n12834), .Y(n3494) );
  OAI21X1 U6696 ( .A(n12747), .B(n12834), .C(n3495), .Y(n7658) );
  NAND2X1 U6697 ( .A(ram[3221]), .B(n12834), .Y(n3495) );
  OAI21X1 U6698 ( .A(n12741), .B(n12834), .C(n3496), .Y(n7659) );
  NAND2X1 U6699 ( .A(ram[3222]), .B(n12834), .Y(n3496) );
  OAI21X1 U6700 ( .A(n12735), .B(n12834), .C(n3497), .Y(n7660) );
  NAND2X1 U6701 ( .A(ram[3223]), .B(n12834), .Y(n3497) );
  OAI21X1 U6702 ( .A(n12729), .B(n12834), .C(n3498), .Y(n7661) );
  NAND2X1 U6703 ( .A(ram[3224]), .B(n12834), .Y(n3498) );
  OAI21X1 U6704 ( .A(n12723), .B(n12834), .C(n3499), .Y(n7662) );
  NAND2X1 U6705 ( .A(ram[3225]), .B(n12834), .Y(n3499) );
  OAI21X1 U6706 ( .A(n12717), .B(n12834), .C(n3500), .Y(n7663) );
  NAND2X1 U6707 ( .A(ram[3226]), .B(n12834), .Y(n3500) );
  OAI21X1 U6708 ( .A(n12711), .B(n12834), .C(n3501), .Y(n7664) );
  NAND2X1 U6709 ( .A(ram[3227]), .B(n12834), .Y(n3501) );
  OAI21X1 U6710 ( .A(n12705), .B(n12834), .C(n3502), .Y(n7665) );
  NAND2X1 U6711 ( .A(ram[3228]), .B(n12834), .Y(n3502) );
  OAI21X1 U6712 ( .A(n12699), .B(n12834), .C(n3503), .Y(n7666) );
  NAND2X1 U6713 ( .A(ram[3229]), .B(n12834), .Y(n3503) );
  OAI21X1 U6714 ( .A(n12693), .B(n12834), .C(n3504), .Y(n7667) );
  NAND2X1 U6715 ( .A(ram[3230]), .B(n12834), .Y(n3504) );
  OAI21X1 U6716 ( .A(n12687), .B(n12834), .C(n3505), .Y(n7668) );
  NAND2X1 U6717 ( .A(ram[3231]), .B(n12834), .Y(n3505) );
  OAI21X1 U6719 ( .A(n12777), .B(n12833), .C(n3507), .Y(n7669) );
  NAND2X1 U6720 ( .A(ram[3232]), .B(n12833), .Y(n3507) );
  OAI21X1 U6721 ( .A(n12771), .B(n12833), .C(n3508), .Y(n7670) );
  NAND2X1 U6722 ( .A(ram[3233]), .B(n12833), .Y(n3508) );
  OAI21X1 U6723 ( .A(n12765), .B(n12833), .C(n3509), .Y(n7671) );
  NAND2X1 U6724 ( .A(ram[3234]), .B(n12833), .Y(n3509) );
  OAI21X1 U6725 ( .A(n12759), .B(n12833), .C(n3510), .Y(n7672) );
  NAND2X1 U6726 ( .A(ram[3235]), .B(n12833), .Y(n3510) );
  OAI21X1 U6727 ( .A(n12753), .B(n12833), .C(n3511), .Y(n7673) );
  NAND2X1 U6728 ( .A(ram[3236]), .B(n12833), .Y(n3511) );
  OAI21X1 U6729 ( .A(n12747), .B(n12833), .C(n3512), .Y(n7674) );
  NAND2X1 U6730 ( .A(ram[3237]), .B(n12833), .Y(n3512) );
  OAI21X1 U6731 ( .A(n12741), .B(n12833), .C(n3513), .Y(n7675) );
  NAND2X1 U6732 ( .A(ram[3238]), .B(n12833), .Y(n3513) );
  OAI21X1 U6733 ( .A(n12735), .B(n12833), .C(n3514), .Y(n7676) );
  NAND2X1 U6734 ( .A(ram[3239]), .B(n12833), .Y(n3514) );
  OAI21X1 U6735 ( .A(n12729), .B(n12833), .C(n3515), .Y(n7677) );
  NAND2X1 U6736 ( .A(ram[3240]), .B(n12833), .Y(n3515) );
  OAI21X1 U6737 ( .A(n12723), .B(n12833), .C(n3516), .Y(n7678) );
  NAND2X1 U6738 ( .A(ram[3241]), .B(n12833), .Y(n3516) );
  OAI21X1 U6739 ( .A(n12717), .B(n12833), .C(n3517), .Y(n7679) );
  NAND2X1 U6740 ( .A(ram[3242]), .B(n12833), .Y(n3517) );
  OAI21X1 U6741 ( .A(n12711), .B(n12833), .C(n3518), .Y(n7680) );
  NAND2X1 U6742 ( .A(ram[3243]), .B(n12833), .Y(n3518) );
  OAI21X1 U6743 ( .A(n12705), .B(n12833), .C(n3519), .Y(n7681) );
  NAND2X1 U6744 ( .A(ram[3244]), .B(n12833), .Y(n3519) );
  OAI21X1 U6745 ( .A(n12699), .B(n12833), .C(n3520), .Y(n7682) );
  NAND2X1 U6746 ( .A(ram[3245]), .B(n12833), .Y(n3520) );
  OAI21X1 U6747 ( .A(n12693), .B(n12833), .C(n3521), .Y(n7683) );
  NAND2X1 U6748 ( .A(ram[3246]), .B(n12833), .Y(n3521) );
  OAI21X1 U6749 ( .A(n12687), .B(n12833), .C(n3522), .Y(n7684) );
  NAND2X1 U6750 ( .A(ram[3247]), .B(n12833), .Y(n3522) );
  OAI21X1 U6752 ( .A(n12777), .B(n12832), .C(n3524), .Y(n7685) );
  NAND2X1 U6753 ( .A(ram[3248]), .B(n12832), .Y(n3524) );
  OAI21X1 U6754 ( .A(n12771), .B(n12832), .C(n3525), .Y(n7686) );
  NAND2X1 U6755 ( .A(ram[3249]), .B(n12832), .Y(n3525) );
  OAI21X1 U6756 ( .A(n12765), .B(n12832), .C(n3526), .Y(n7687) );
  NAND2X1 U6757 ( .A(ram[3250]), .B(n12832), .Y(n3526) );
  OAI21X1 U6758 ( .A(n12759), .B(n12832), .C(n3527), .Y(n7688) );
  NAND2X1 U6759 ( .A(ram[3251]), .B(n12832), .Y(n3527) );
  OAI21X1 U6760 ( .A(n12753), .B(n12832), .C(n3528), .Y(n7689) );
  NAND2X1 U6761 ( .A(ram[3252]), .B(n12832), .Y(n3528) );
  OAI21X1 U6762 ( .A(n12747), .B(n12832), .C(n3529), .Y(n7690) );
  NAND2X1 U6763 ( .A(ram[3253]), .B(n12832), .Y(n3529) );
  OAI21X1 U6764 ( .A(n12741), .B(n12832), .C(n3530), .Y(n7691) );
  NAND2X1 U6765 ( .A(ram[3254]), .B(n12832), .Y(n3530) );
  OAI21X1 U6766 ( .A(n12735), .B(n12832), .C(n3531), .Y(n7692) );
  NAND2X1 U6767 ( .A(ram[3255]), .B(n12832), .Y(n3531) );
  OAI21X1 U6768 ( .A(n12729), .B(n12832), .C(n3532), .Y(n7693) );
  NAND2X1 U6769 ( .A(ram[3256]), .B(n12832), .Y(n3532) );
  OAI21X1 U6770 ( .A(n12723), .B(n12832), .C(n3533), .Y(n7694) );
  NAND2X1 U6771 ( .A(ram[3257]), .B(n12832), .Y(n3533) );
  OAI21X1 U6772 ( .A(n12717), .B(n12832), .C(n3534), .Y(n7695) );
  NAND2X1 U6773 ( .A(ram[3258]), .B(n12832), .Y(n3534) );
  OAI21X1 U6774 ( .A(n12711), .B(n12832), .C(n3535), .Y(n7696) );
  NAND2X1 U6775 ( .A(ram[3259]), .B(n12832), .Y(n3535) );
  OAI21X1 U6776 ( .A(n12705), .B(n12832), .C(n3536), .Y(n7697) );
  NAND2X1 U6777 ( .A(ram[3260]), .B(n12832), .Y(n3536) );
  OAI21X1 U6778 ( .A(n12699), .B(n12832), .C(n3537), .Y(n7698) );
  NAND2X1 U6779 ( .A(ram[3261]), .B(n12832), .Y(n3537) );
  OAI21X1 U6780 ( .A(n12693), .B(n12832), .C(n3538), .Y(n7699) );
  NAND2X1 U6781 ( .A(ram[3262]), .B(n12832), .Y(n3538) );
  OAI21X1 U6782 ( .A(n12687), .B(n12832), .C(n3539), .Y(n7700) );
  NAND2X1 U6783 ( .A(ram[3263]), .B(n12832), .Y(n3539) );
  OAI21X1 U6785 ( .A(n12777), .B(n12831), .C(n3541), .Y(n7701) );
  NAND2X1 U6786 ( .A(ram[3264]), .B(n12831), .Y(n3541) );
  OAI21X1 U6787 ( .A(n12771), .B(n12831), .C(n3542), .Y(n7702) );
  NAND2X1 U6788 ( .A(ram[3265]), .B(n12831), .Y(n3542) );
  OAI21X1 U6789 ( .A(n12765), .B(n12831), .C(n3543), .Y(n7703) );
  NAND2X1 U6790 ( .A(ram[3266]), .B(n12831), .Y(n3543) );
  OAI21X1 U6791 ( .A(n12759), .B(n12831), .C(n3544), .Y(n7704) );
  NAND2X1 U6792 ( .A(ram[3267]), .B(n12831), .Y(n3544) );
  OAI21X1 U6793 ( .A(n12753), .B(n12831), .C(n3545), .Y(n7705) );
  NAND2X1 U6794 ( .A(ram[3268]), .B(n12831), .Y(n3545) );
  OAI21X1 U6795 ( .A(n12747), .B(n12831), .C(n3546), .Y(n7706) );
  NAND2X1 U6796 ( .A(ram[3269]), .B(n12831), .Y(n3546) );
  OAI21X1 U6797 ( .A(n12741), .B(n12831), .C(n3547), .Y(n7707) );
  NAND2X1 U6798 ( .A(ram[3270]), .B(n12831), .Y(n3547) );
  OAI21X1 U6799 ( .A(n12735), .B(n12831), .C(n3548), .Y(n7708) );
  NAND2X1 U6800 ( .A(ram[3271]), .B(n12831), .Y(n3548) );
  OAI21X1 U6801 ( .A(n12729), .B(n12831), .C(n3549), .Y(n7709) );
  NAND2X1 U6802 ( .A(ram[3272]), .B(n12831), .Y(n3549) );
  OAI21X1 U6803 ( .A(n12723), .B(n12831), .C(n3550), .Y(n7710) );
  NAND2X1 U6804 ( .A(ram[3273]), .B(n12831), .Y(n3550) );
  OAI21X1 U6805 ( .A(n12717), .B(n12831), .C(n3551), .Y(n7711) );
  NAND2X1 U6806 ( .A(ram[3274]), .B(n12831), .Y(n3551) );
  OAI21X1 U6807 ( .A(n12711), .B(n12831), .C(n3552), .Y(n7712) );
  NAND2X1 U6808 ( .A(ram[3275]), .B(n12831), .Y(n3552) );
  OAI21X1 U6809 ( .A(n12705), .B(n12831), .C(n3553), .Y(n7713) );
  NAND2X1 U6810 ( .A(ram[3276]), .B(n12831), .Y(n3553) );
  OAI21X1 U6811 ( .A(n12699), .B(n12831), .C(n3554), .Y(n7714) );
  NAND2X1 U6812 ( .A(ram[3277]), .B(n12831), .Y(n3554) );
  OAI21X1 U6813 ( .A(n12693), .B(n12831), .C(n3555), .Y(n7715) );
  NAND2X1 U6814 ( .A(ram[3278]), .B(n12831), .Y(n3555) );
  OAI21X1 U6815 ( .A(n12687), .B(n12831), .C(n3556), .Y(n7716) );
  NAND2X1 U6816 ( .A(ram[3279]), .B(n12831), .Y(n3556) );
  OAI21X1 U6818 ( .A(n12777), .B(n12830), .C(n3558), .Y(n7717) );
  NAND2X1 U6819 ( .A(ram[3280]), .B(n12830), .Y(n3558) );
  OAI21X1 U6820 ( .A(n12771), .B(n12830), .C(n3559), .Y(n7718) );
  NAND2X1 U6821 ( .A(ram[3281]), .B(n12830), .Y(n3559) );
  OAI21X1 U6822 ( .A(n12765), .B(n12830), .C(n3560), .Y(n7719) );
  NAND2X1 U6823 ( .A(ram[3282]), .B(n12830), .Y(n3560) );
  OAI21X1 U6824 ( .A(n12759), .B(n12830), .C(n3561), .Y(n7720) );
  NAND2X1 U6825 ( .A(ram[3283]), .B(n12830), .Y(n3561) );
  OAI21X1 U6826 ( .A(n12753), .B(n12830), .C(n3562), .Y(n7721) );
  NAND2X1 U6827 ( .A(ram[3284]), .B(n12830), .Y(n3562) );
  OAI21X1 U6828 ( .A(n12747), .B(n12830), .C(n3563), .Y(n7722) );
  NAND2X1 U6829 ( .A(ram[3285]), .B(n12830), .Y(n3563) );
  OAI21X1 U6830 ( .A(n12741), .B(n12830), .C(n3564), .Y(n7723) );
  NAND2X1 U6831 ( .A(ram[3286]), .B(n12830), .Y(n3564) );
  OAI21X1 U6832 ( .A(n12735), .B(n12830), .C(n3565), .Y(n7724) );
  NAND2X1 U6833 ( .A(ram[3287]), .B(n12830), .Y(n3565) );
  OAI21X1 U6834 ( .A(n12729), .B(n12830), .C(n3566), .Y(n7725) );
  NAND2X1 U6835 ( .A(ram[3288]), .B(n12830), .Y(n3566) );
  OAI21X1 U6836 ( .A(n12723), .B(n12830), .C(n3567), .Y(n7726) );
  NAND2X1 U6837 ( .A(ram[3289]), .B(n12830), .Y(n3567) );
  OAI21X1 U6838 ( .A(n12717), .B(n12830), .C(n3568), .Y(n7727) );
  NAND2X1 U6839 ( .A(ram[3290]), .B(n12830), .Y(n3568) );
  OAI21X1 U6840 ( .A(n12711), .B(n12830), .C(n3569), .Y(n7728) );
  NAND2X1 U6841 ( .A(ram[3291]), .B(n12830), .Y(n3569) );
  OAI21X1 U6842 ( .A(n12705), .B(n12830), .C(n3570), .Y(n7729) );
  NAND2X1 U6843 ( .A(ram[3292]), .B(n12830), .Y(n3570) );
  OAI21X1 U6844 ( .A(n12699), .B(n12830), .C(n3571), .Y(n7730) );
  NAND2X1 U6845 ( .A(ram[3293]), .B(n12830), .Y(n3571) );
  OAI21X1 U6846 ( .A(n12693), .B(n12830), .C(n3572), .Y(n7731) );
  NAND2X1 U6847 ( .A(ram[3294]), .B(n12830), .Y(n3572) );
  OAI21X1 U6848 ( .A(n12687), .B(n12830), .C(n3573), .Y(n7732) );
  NAND2X1 U6849 ( .A(ram[3295]), .B(n12830), .Y(n3573) );
  OAI21X1 U6851 ( .A(n12777), .B(n12829), .C(n3575), .Y(n7733) );
  NAND2X1 U6852 ( .A(ram[3296]), .B(n12829), .Y(n3575) );
  OAI21X1 U6853 ( .A(n12771), .B(n12829), .C(n3576), .Y(n7734) );
  NAND2X1 U6854 ( .A(ram[3297]), .B(n12829), .Y(n3576) );
  OAI21X1 U6855 ( .A(n12765), .B(n12829), .C(n3577), .Y(n7735) );
  NAND2X1 U6856 ( .A(ram[3298]), .B(n12829), .Y(n3577) );
  OAI21X1 U6857 ( .A(n12759), .B(n12829), .C(n3578), .Y(n7736) );
  NAND2X1 U6858 ( .A(ram[3299]), .B(n12829), .Y(n3578) );
  OAI21X1 U6859 ( .A(n12753), .B(n12829), .C(n3579), .Y(n7737) );
  NAND2X1 U6860 ( .A(ram[3300]), .B(n12829), .Y(n3579) );
  OAI21X1 U6861 ( .A(n12747), .B(n12829), .C(n3580), .Y(n7738) );
  NAND2X1 U6862 ( .A(ram[3301]), .B(n12829), .Y(n3580) );
  OAI21X1 U6863 ( .A(n12741), .B(n12829), .C(n3581), .Y(n7739) );
  NAND2X1 U6864 ( .A(ram[3302]), .B(n12829), .Y(n3581) );
  OAI21X1 U6865 ( .A(n12735), .B(n12829), .C(n3582), .Y(n7740) );
  NAND2X1 U6866 ( .A(ram[3303]), .B(n12829), .Y(n3582) );
  OAI21X1 U6867 ( .A(n12729), .B(n12829), .C(n3583), .Y(n7741) );
  NAND2X1 U6868 ( .A(ram[3304]), .B(n12829), .Y(n3583) );
  OAI21X1 U6869 ( .A(n12723), .B(n12829), .C(n3584), .Y(n7742) );
  NAND2X1 U6870 ( .A(ram[3305]), .B(n12829), .Y(n3584) );
  OAI21X1 U6871 ( .A(n12717), .B(n12829), .C(n3585), .Y(n7743) );
  NAND2X1 U6872 ( .A(ram[3306]), .B(n12829), .Y(n3585) );
  OAI21X1 U6873 ( .A(n12711), .B(n12829), .C(n3586), .Y(n7744) );
  NAND2X1 U6874 ( .A(ram[3307]), .B(n12829), .Y(n3586) );
  OAI21X1 U6875 ( .A(n12705), .B(n12829), .C(n3587), .Y(n7745) );
  NAND2X1 U6876 ( .A(ram[3308]), .B(n12829), .Y(n3587) );
  OAI21X1 U6877 ( .A(n12699), .B(n12829), .C(n3588), .Y(n7746) );
  NAND2X1 U6878 ( .A(ram[3309]), .B(n12829), .Y(n3588) );
  OAI21X1 U6879 ( .A(n12693), .B(n12829), .C(n3589), .Y(n7747) );
  NAND2X1 U6880 ( .A(ram[3310]), .B(n12829), .Y(n3589) );
  OAI21X1 U6881 ( .A(n12687), .B(n12829), .C(n3590), .Y(n7748) );
  NAND2X1 U6882 ( .A(ram[3311]), .B(n12829), .Y(n3590) );
  OAI21X1 U6884 ( .A(n12777), .B(n12828), .C(n3592), .Y(n7749) );
  NAND2X1 U6885 ( .A(ram[3312]), .B(n12828), .Y(n3592) );
  OAI21X1 U6886 ( .A(n12771), .B(n12828), .C(n3593), .Y(n7750) );
  NAND2X1 U6887 ( .A(ram[3313]), .B(n12828), .Y(n3593) );
  OAI21X1 U6888 ( .A(n12765), .B(n12828), .C(n3594), .Y(n7751) );
  NAND2X1 U6889 ( .A(ram[3314]), .B(n12828), .Y(n3594) );
  OAI21X1 U6890 ( .A(n12759), .B(n12828), .C(n3595), .Y(n7752) );
  NAND2X1 U6891 ( .A(ram[3315]), .B(n12828), .Y(n3595) );
  OAI21X1 U6892 ( .A(n12753), .B(n12828), .C(n3596), .Y(n7753) );
  NAND2X1 U6893 ( .A(ram[3316]), .B(n12828), .Y(n3596) );
  OAI21X1 U6894 ( .A(n12747), .B(n12828), .C(n3597), .Y(n7754) );
  NAND2X1 U6895 ( .A(ram[3317]), .B(n12828), .Y(n3597) );
  OAI21X1 U6896 ( .A(n12741), .B(n12828), .C(n3598), .Y(n7755) );
  NAND2X1 U6897 ( .A(ram[3318]), .B(n12828), .Y(n3598) );
  OAI21X1 U6898 ( .A(n12735), .B(n12828), .C(n3599), .Y(n7756) );
  NAND2X1 U6899 ( .A(ram[3319]), .B(n12828), .Y(n3599) );
  OAI21X1 U6900 ( .A(n12729), .B(n12828), .C(n3600), .Y(n7757) );
  NAND2X1 U6901 ( .A(ram[3320]), .B(n12828), .Y(n3600) );
  OAI21X1 U6902 ( .A(n12723), .B(n12828), .C(n3601), .Y(n7758) );
  NAND2X1 U6903 ( .A(ram[3321]), .B(n12828), .Y(n3601) );
  OAI21X1 U6904 ( .A(n12717), .B(n12828), .C(n3602), .Y(n7759) );
  NAND2X1 U6905 ( .A(ram[3322]), .B(n12828), .Y(n3602) );
  OAI21X1 U6906 ( .A(n12711), .B(n12828), .C(n3603), .Y(n7760) );
  NAND2X1 U6907 ( .A(ram[3323]), .B(n12828), .Y(n3603) );
  OAI21X1 U6908 ( .A(n12705), .B(n12828), .C(n3604), .Y(n7761) );
  NAND2X1 U6909 ( .A(ram[3324]), .B(n12828), .Y(n3604) );
  OAI21X1 U6910 ( .A(n12699), .B(n12828), .C(n3605), .Y(n7762) );
  NAND2X1 U6911 ( .A(ram[3325]), .B(n12828), .Y(n3605) );
  OAI21X1 U6912 ( .A(n12693), .B(n12828), .C(n3606), .Y(n7763) );
  NAND2X1 U6913 ( .A(ram[3326]), .B(n12828), .Y(n3606) );
  OAI21X1 U6914 ( .A(n12687), .B(n12828), .C(n3607), .Y(n7764) );
  NAND2X1 U6915 ( .A(ram[3327]), .B(n12828), .Y(n3607) );
  NAND3X1 U6917 ( .A(mem_write_en), .B(n327), .C(n3609), .Y(n3608) );
  NOR2X1 U6918 ( .A(mem_access_addr[4]), .B(mem_access_addr[5]), .Y(n327) );
  OAI21X1 U6919 ( .A(n12778), .B(n12827), .C(n3611), .Y(n7765) );
  NAND2X1 U6920 ( .A(ram[3328]), .B(n12827), .Y(n3611) );
  OAI21X1 U6921 ( .A(n12772), .B(n12827), .C(n3612), .Y(n7766) );
  NAND2X1 U6922 ( .A(ram[3329]), .B(n12827), .Y(n3612) );
  OAI21X1 U6923 ( .A(n12766), .B(n12827), .C(n3613), .Y(n7767) );
  NAND2X1 U6924 ( .A(ram[3330]), .B(n12827), .Y(n3613) );
  OAI21X1 U6925 ( .A(n12760), .B(n12827), .C(n3614), .Y(n7768) );
  NAND2X1 U6926 ( .A(ram[3331]), .B(n12827), .Y(n3614) );
  OAI21X1 U6927 ( .A(n12754), .B(n12827), .C(n3615), .Y(n7769) );
  NAND2X1 U6928 ( .A(ram[3332]), .B(n12827), .Y(n3615) );
  OAI21X1 U6929 ( .A(n12748), .B(n12827), .C(n3616), .Y(n7770) );
  NAND2X1 U6930 ( .A(ram[3333]), .B(n12827), .Y(n3616) );
  OAI21X1 U6931 ( .A(n12742), .B(n12827), .C(n3617), .Y(n7771) );
  NAND2X1 U6932 ( .A(ram[3334]), .B(n12827), .Y(n3617) );
  OAI21X1 U6933 ( .A(n12736), .B(n12827), .C(n3618), .Y(n7772) );
  NAND2X1 U6934 ( .A(ram[3335]), .B(n12827), .Y(n3618) );
  OAI21X1 U6935 ( .A(n12730), .B(n12827), .C(n3619), .Y(n7773) );
  NAND2X1 U6936 ( .A(ram[3336]), .B(n12827), .Y(n3619) );
  OAI21X1 U6937 ( .A(n12724), .B(n12827), .C(n3620), .Y(n7774) );
  NAND2X1 U6938 ( .A(ram[3337]), .B(n12827), .Y(n3620) );
  OAI21X1 U6939 ( .A(n12718), .B(n12827), .C(n3621), .Y(n7775) );
  NAND2X1 U6940 ( .A(ram[3338]), .B(n12827), .Y(n3621) );
  OAI21X1 U6941 ( .A(n12712), .B(n12827), .C(n3622), .Y(n7776) );
  NAND2X1 U6942 ( .A(ram[3339]), .B(n12827), .Y(n3622) );
  OAI21X1 U6943 ( .A(n12706), .B(n12827), .C(n3623), .Y(n7777) );
  NAND2X1 U6944 ( .A(ram[3340]), .B(n12827), .Y(n3623) );
  OAI21X1 U6945 ( .A(n12700), .B(n12827), .C(n3624), .Y(n7778) );
  NAND2X1 U6946 ( .A(ram[3341]), .B(n12827), .Y(n3624) );
  OAI21X1 U6947 ( .A(n12694), .B(n12827), .C(n3625), .Y(n7779) );
  NAND2X1 U6948 ( .A(ram[3342]), .B(n12827), .Y(n3625) );
  OAI21X1 U6949 ( .A(n12688), .B(n12827), .C(n3626), .Y(n7780) );
  NAND2X1 U6950 ( .A(ram[3343]), .B(n12827), .Y(n3626) );
  OAI21X1 U6952 ( .A(n12778), .B(n12826), .C(n3628), .Y(n7781) );
  NAND2X1 U6953 ( .A(ram[3344]), .B(n12826), .Y(n3628) );
  OAI21X1 U6954 ( .A(n12772), .B(n12826), .C(n3629), .Y(n7782) );
  NAND2X1 U6955 ( .A(ram[3345]), .B(n12826), .Y(n3629) );
  OAI21X1 U6956 ( .A(n12766), .B(n12826), .C(n3630), .Y(n7783) );
  NAND2X1 U6957 ( .A(ram[3346]), .B(n12826), .Y(n3630) );
  OAI21X1 U6958 ( .A(n12760), .B(n12826), .C(n3631), .Y(n7784) );
  NAND2X1 U6959 ( .A(ram[3347]), .B(n12826), .Y(n3631) );
  OAI21X1 U6960 ( .A(n12754), .B(n12826), .C(n3632), .Y(n7785) );
  NAND2X1 U6961 ( .A(ram[3348]), .B(n12826), .Y(n3632) );
  OAI21X1 U6962 ( .A(n12748), .B(n12826), .C(n3633), .Y(n7786) );
  NAND2X1 U6963 ( .A(ram[3349]), .B(n12826), .Y(n3633) );
  OAI21X1 U6964 ( .A(n12742), .B(n12826), .C(n3634), .Y(n7787) );
  NAND2X1 U6965 ( .A(ram[3350]), .B(n12826), .Y(n3634) );
  OAI21X1 U6966 ( .A(n12736), .B(n12826), .C(n3635), .Y(n7788) );
  NAND2X1 U6967 ( .A(ram[3351]), .B(n12826), .Y(n3635) );
  OAI21X1 U6968 ( .A(n12730), .B(n12826), .C(n3636), .Y(n7789) );
  NAND2X1 U6969 ( .A(ram[3352]), .B(n12826), .Y(n3636) );
  OAI21X1 U6970 ( .A(n12724), .B(n12826), .C(n3637), .Y(n7790) );
  NAND2X1 U6971 ( .A(ram[3353]), .B(n12826), .Y(n3637) );
  OAI21X1 U6972 ( .A(n12718), .B(n12826), .C(n3638), .Y(n7791) );
  NAND2X1 U6973 ( .A(ram[3354]), .B(n12826), .Y(n3638) );
  OAI21X1 U6974 ( .A(n12712), .B(n12826), .C(n3639), .Y(n7792) );
  NAND2X1 U6975 ( .A(ram[3355]), .B(n12826), .Y(n3639) );
  OAI21X1 U6976 ( .A(n12706), .B(n12826), .C(n3640), .Y(n7793) );
  NAND2X1 U6977 ( .A(ram[3356]), .B(n12826), .Y(n3640) );
  OAI21X1 U6978 ( .A(n12700), .B(n12826), .C(n3641), .Y(n7794) );
  NAND2X1 U6979 ( .A(ram[3357]), .B(n12826), .Y(n3641) );
  OAI21X1 U6980 ( .A(n12694), .B(n12826), .C(n3642), .Y(n7795) );
  NAND2X1 U6981 ( .A(ram[3358]), .B(n12826), .Y(n3642) );
  OAI21X1 U6982 ( .A(n12688), .B(n12826), .C(n3643), .Y(n7796) );
  NAND2X1 U6983 ( .A(ram[3359]), .B(n12826), .Y(n3643) );
  OAI21X1 U6985 ( .A(n12778), .B(n12825), .C(n3645), .Y(n7797) );
  NAND2X1 U6986 ( .A(ram[3360]), .B(n12825), .Y(n3645) );
  OAI21X1 U6987 ( .A(n12772), .B(n12825), .C(n3646), .Y(n7798) );
  NAND2X1 U6988 ( .A(ram[3361]), .B(n12825), .Y(n3646) );
  OAI21X1 U6989 ( .A(n12766), .B(n12825), .C(n3647), .Y(n7799) );
  NAND2X1 U6990 ( .A(ram[3362]), .B(n12825), .Y(n3647) );
  OAI21X1 U6991 ( .A(n12760), .B(n12825), .C(n3648), .Y(n7800) );
  NAND2X1 U6992 ( .A(ram[3363]), .B(n12825), .Y(n3648) );
  OAI21X1 U6993 ( .A(n12754), .B(n12825), .C(n3649), .Y(n7801) );
  NAND2X1 U6994 ( .A(ram[3364]), .B(n12825), .Y(n3649) );
  OAI21X1 U6995 ( .A(n12748), .B(n12825), .C(n3650), .Y(n7802) );
  NAND2X1 U6996 ( .A(ram[3365]), .B(n12825), .Y(n3650) );
  OAI21X1 U6997 ( .A(n12742), .B(n12825), .C(n3651), .Y(n7803) );
  NAND2X1 U6998 ( .A(ram[3366]), .B(n12825), .Y(n3651) );
  OAI21X1 U6999 ( .A(n12736), .B(n12825), .C(n3652), .Y(n7804) );
  NAND2X1 U7000 ( .A(ram[3367]), .B(n12825), .Y(n3652) );
  OAI21X1 U7001 ( .A(n12730), .B(n12825), .C(n3653), .Y(n7805) );
  NAND2X1 U7002 ( .A(ram[3368]), .B(n12825), .Y(n3653) );
  OAI21X1 U7003 ( .A(n12724), .B(n12825), .C(n3654), .Y(n7806) );
  NAND2X1 U7004 ( .A(ram[3369]), .B(n12825), .Y(n3654) );
  OAI21X1 U7005 ( .A(n12718), .B(n12825), .C(n3655), .Y(n7807) );
  NAND2X1 U7006 ( .A(ram[3370]), .B(n12825), .Y(n3655) );
  OAI21X1 U7007 ( .A(n12712), .B(n12825), .C(n3656), .Y(n7808) );
  NAND2X1 U7008 ( .A(ram[3371]), .B(n12825), .Y(n3656) );
  OAI21X1 U7009 ( .A(n12706), .B(n12825), .C(n3657), .Y(n7809) );
  NAND2X1 U7010 ( .A(ram[3372]), .B(n12825), .Y(n3657) );
  OAI21X1 U7011 ( .A(n12700), .B(n12825), .C(n3658), .Y(n7810) );
  NAND2X1 U7012 ( .A(ram[3373]), .B(n12825), .Y(n3658) );
  OAI21X1 U7013 ( .A(n12694), .B(n12825), .C(n3659), .Y(n7811) );
  NAND2X1 U7014 ( .A(ram[3374]), .B(n12825), .Y(n3659) );
  OAI21X1 U7015 ( .A(n12688), .B(n12825), .C(n3660), .Y(n7812) );
  NAND2X1 U7016 ( .A(ram[3375]), .B(n12825), .Y(n3660) );
  OAI21X1 U7018 ( .A(n12778), .B(n12824), .C(n3662), .Y(n7813) );
  NAND2X1 U7019 ( .A(ram[3376]), .B(n12824), .Y(n3662) );
  OAI21X1 U7020 ( .A(n12772), .B(n12824), .C(n3663), .Y(n7814) );
  NAND2X1 U7021 ( .A(ram[3377]), .B(n12824), .Y(n3663) );
  OAI21X1 U7022 ( .A(n12766), .B(n12824), .C(n3664), .Y(n7815) );
  NAND2X1 U7023 ( .A(ram[3378]), .B(n12824), .Y(n3664) );
  OAI21X1 U7024 ( .A(n12760), .B(n12824), .C(n3665), .Y(n7816) );
  NAND2X1 U7025 ( .A(ram[3379]), .B(n12824), .Y(n3665) );
  OAI21X1 U7026 ( .A(n12754), .B(n12824), .C(n3666), .Y(n7817) );
  NAND2X1 U7027 ( .A(ram[3380]), .B(n12824), .Y(n3666) );
  OAI21X1 U7028 ( .A(n12748), .B(n12824), .C(n3667), .Y(n7818) );
  NAND2X1 U7029 ( .A(ram[3381]), .B(n12824), .Y(n3667) );
  OAI21X1 U7030 ( .A(n12742), .B(n12824), .C(n3668), .Y(n7819) );
  NAND2X1 U7031 ( .A(ram[3382]), .B(n12824), .Y(n3668) );
  OAI21X1 U7032 ( .A(n12736), .B(n12824), .C(n3669), .Y(n7820) );
  NAND2X1 U7033 ( .A(ram[3383]), .B(n12824), .Y(n3669) );
  OAI21X1 U7034 ( .A(n12730), .B(n12824), .C(n3670), .Y(n7821) );
  NAND2X1 U7035 ( .A(ram[3384]), .B(n12824), .Y(n3670) );
  OAI21X1 U7036 ( .A(n12724), .B(n12824), .C(n3671), .Y(n7822) );
  NAND2X1 U7037 ( .A(ram[3385]), .B(n12824), .Y(n3671) );
  OAI21X1 U7038 ( .A(n12718), .B(n12824), .C(n3672), .Y(n7823) );
  NAND2X1 U7039 ( .A(ram[3386]), .B(n12824), .Y(n3672) );
  OAI21X1 U7040 ( .A(n12712), .B(n12824), .C(n3673), .Y(n7824) );
  NAND2X1 U7041 ( .A(ram[3387]), .B(n12824), .Y(n3673) );
  OAI21X1 U7042 ( .A(n12706), .B(n12824), .C(n3674), .Y(n7825) );
  NAND2X1 U7043 ( .A(ram[3388]), .B(n12824), .Y(n3674) );
  OAI21X1 U7044 ( .A(n12700), .B(n12824), .C(n3675), .Y(n7826) );
  NAND2X1 U7045 ( .A(ram[3389]), .B(n12824), .Y(n3675) );
  OAI21X1 U7046 ( .A(n12694), .B(n12824), .C(n3676), .Y(n7827) );
  NAND2X1 U7047 ( .A(ram[3390]), .B(n12824), .Y(n3676) );
  OAI21X1 U7048 ( .A(n12688), .B(n12824), .C(n3677), .Y(n7828) );
  NAND2X1 U7049 ( .A(ram[3391]), .B(n12824), .Y(n3677) );
  OAI21X1 U7051 ( .A(n12778), .B(n12823), .C(n3679), .Y(n7829) );
  NAND2X1 U7052 ( .A(ram[3392]), .B(n12823), .Y(n3679) );
  OAI21X1 U7053 ( .A(n12772), .B(n12823), .C(n3680), .Y(n7830) );
  NAND2X1 U7054 ( .A(ram[3393]), .B(n12823), .Y(n3680) );
  OAI21X1 U7055 ( .A(n12766), .B(n12823), .C(n3681), .Y(n7831) );
  NAND2X1 U7056 ( .A(ram[3394]), .B(n12823), .Y(n3681) );
  OAI21X1 U7057 ( .A(n12760), .B(n12823), .C(n3682), .Y(n7832) );
  NAND2X1 U7058 ( .A(ram[3395]), .B(n12823), .Y(n3682) );
  OAI21X1 U7059 ( .A(n12754), .B(n12823), .C(n3683), .Y(n7833) );
  NAND2X1 U7060 ( .A(ram[3396]), .B(n12823), .Y(n3683) );
  OAI21X1 U7061 ( .A(n12748), .B(n12823), .C(n3684), .Y(n7834) );
  NAND2X1 U7062 ( .A(ram[3397]), .B(n12823), .Y(n3684) );
  OAI21X1 U7063 ( .A(n12742), .B(n12823), .C(n3685), .Y(n7835) );
  NAND2X1 U7064 ( .A(ram[3398]), .B(n12823), .Y(n3685) );
  OAI21X1 U7065 ( .A(n12736), .B(n12823), .C(n3686), .Y(n7836) );
  NAND2X1 U7066 ( .A(ram[3399]), .B(n12823), .Y(n3686) );
  OAI21X1 U7067 ( .A(n12730), .B(n12823), .C(n3687), .Y(n7837) );
  NAND2X1 U7068 ( .A(ram[3400]), .B(n12823), .Y(n3687) );
  OAI21X1 U7069 ( .A(n12724), .B(n12823), .C(n3688), .Y(n7838) );
  NAND2X1 U7070 ( .A(ram[3401]), .B(n12823), .Y(n3688) );
  OAI21X1 U7071 ( .A(n12718), .B(n12823), .C(n3689), .Y(n7839) );
  NAND2X1 U7072 ( .A(ram[3402]), .B(n12823), .Y(n3689) );
  OAI21X1 U7073 ( .A(n12712), .B(n12823), .C(n3690), .Y(n7840) );
  NAND2X1 U7074 ( .A(ram[3403]), .B(n12823), .Y(n3690) );
  OAI21X1 U7075 ( .A(n12706), .B(n12823), .C(n3691), .Y(n7841) );
  NAND2X1 U7076 ( .A(ram[3404]), .B(n12823), .Y(n3691) );
  OAI21X1 U7077 ( .A(n12700), .B(n12823), .C(n3692), .Y(n7842) );
  NAND2X1 U7078 ( .A(ram[3405]), .B(n12823), .Y(n3692) );
  OAI21X1 U7079 ( .A(n12694), .B(n12823), .C(n3693), .Y(n7843) );
  NAND2X1 U7080 ( .A(ram[3406]), .B(n12823), .Y(n3693) );
  OAI21X1 U7081 ( .A(n12688), .B(n12823), .C(n3694), .Y(n7844) );
  NAND2X1 U7082 ( .A(ram[3407]), .B(n12823), .Y(n3694) );
  OAI21X1 U7084 ( .A(n12778), .B(n12822), .C(n3696), .Y(n7845) );
  NAND2X1 U7085 ( .A(ram[3408]), .B(n12822), .Y(n3696) );
  OAI21X1 U7086 ( .A(n12772), .B(n12822), .C(n3697), .Y(n7846) );
  NAND2X1 U7087 ( .A(ram[3409]), .B(n12822), .Y(n3697) );
  OAI21X1 U7088 ( .A(n12766), .B(n12822), .C(n3698), .Y(n7847) );
  NAND2X1 U7089 ( .A(ram[3410]), .B(n12822), .Y(n3698) );
  OAI21X1 U7090 ( .A(n12760), .B(n12822), .C(n3699), .Y(n7848) );
  NAND2X1 U7091 ( .A(ram[3411]), .B(n12822), .Y(n3699) );
  OAI21X1 U7092 ( .A(n12754), .B(n12822), .C(n3700), .Y(n7849) );
  NAND2X1 U7093 ( .A(ram[3412]), .B(n12822), .Y(n3700) );
  OAI21X1 U7094 ( .A(n12748), .B(n12822), .C(n3701), .Y(n7850) );
  NAND2X1 U7095 ( .A(ram[3413]), .B(n12822), .Y(n3701) );
  OAI21X1 U7096 ( .A(n12742), .B(n12822), .C(n3702), .Y(n7851) );
  NAND2X1 U7097 ( .A(ram[3414]), .B(n12822), .Y(n3702) );
  OAI21X1 U7098 ( .A(n12736), .B(n12822), .C(n3703), .Y(n7852) );
  NAND2X1 U7099 ( .A(ram[3415]), .B(n12822), .Y(n3703) );
  OAI21X1 U7100 ( .A(n12730), .B(n12822), .C(n3704), .Y(n7853) );
  NAND2X1 U7101 ( .A(ram[3416]), .B(n12822), .Y(n3704) );
  OAI21X1 U7102 ( .A(n12724), .B(n12822), .C(n3705), .Y(n7854) );
  NAND2X1 U7103 ( .A(ram[3417]), .B(n12822), .Y(n3705) );
  OAI21X1 U7104 ( .A(n12718), .B(n12822), .C(n3706), .Y(n7855) );
  NAND2X1 U7105 ( .A(ram[3418]), .B(n12822), .Y(n3706) );
  OAI21X1 U7106 ( .A(n12712), .B(n12822), .C(n3707), .Y(n7856) );
  NAND2X1 U7107 ( .A(ram[3419]), .B(n12822), .Y(n3707) );
  OAI21X1 U7108 ( .A(n12706), .B(n12822), .C(n3708), .Y(n7857) );
  NAND2X1 U7109 ( .A(ram[3420]), .B(n12822), .Y(n3708) );
  OAI21X1 U7110 ( .A(n12700), .B(n12822), .C(n3709), .Y(n7858) );
  NAND2X1 U7111 ( .A(ram[3421]), .B(n12822), .Y(n3709) );
  OAI21X1 U7112 ( .A(n12694), .B(n12822), .C(n3710), .Y(n7859) );
  NAND2X1 U7113 ( .A(ram[3422]), .B(n12822), .Y(n3710) );
  OAI21X1 U7114 ( .A(n12688), .B(n12822), .C(n3711), .Y(n7860) );
  NAND2X1 U7115 ( .A(ram[3423]), .B(n12822), .Y(n3711) );
  OAI21X1 U7117 ( .A(n12778), .B(n12821), .C(n3713), .Y(n7861) );
  NAND2X1 U7118 ( .A(ram[3424]), .B(n12821), .Y(n3713) );
  OAI21X1 U7119 ( .A(n12772), .B(n12821), .C(n3714), .Y(n7862) );
  NAND2X1 U7120 ( .A(ram[3425]), .B(n12821), .Y(n3714) );
  OAI21X1 U7121 ( .A(n12766), .B(n12821), .C(n3715), .Y(n7863) );
  NAND2X1 U7122 ( .A(ram[3426]), .B(n12821), .Y(n3715) );
  OAI21X1 U7123 ( .A(n12760), .B(n12821), .C(n3716), .Y(n7864) );
  NAND2X1 U7124 ( .A(ram[3427]), .B(n12821), .Y(n3716) );
  OAI21X1 U7125 ( .A(n12754), .B(n12821), .C(n3717), .Y(n7865) );
  NAND2X1 U7126 ( .A(ram[3428]), .B(n12821), .Y(n3717) );
  OAI21X1 U7127 ( .A(n12748), .B(n12821), .C(n3718), .Y(n7866) );
  NAND2X1 U7128 ( .A(ram[3429]), .B(n12821), .Y(n3718) );
  OAI21X1 U7129 ( .A(n12742), .B(n12821), .C(n3719), .Y(n7867) );
  NAND2X1 U7130 ( .A(ram[3430]), .B(n12821), .Y(n3719) );
  OAI21X1 U7131 ( .A(n12736), .B(n12821), .C(n3720), .Y(n7868) );
  NAND2X1 U7132 ( .A(ram[3431]), .B(n12821), .Y(n3720) );
  OAI21X1 U7133 ( .A(n12730), .B(n12821), .C(n3721), .Y(n7869) );
  NAND2X1 U7134 ( .A(ram[3432]), .B(n12821), .Y(n3721) );
  OAI21X1 U7135 ( .A(n12724), .B(n12821), .C(n3722), .Y(n7870) );
  NAND2X1 U7136 ( .A(ram[3433]), .B(n12821), .Y(n3722) );
  OAI21X1 U7137 ( .A(n12718), .B(n12821), .C(n3723), .Y(n7871) );
  NAND2X1 U7138 ( .A(ram[3434]), .B(n12821), .Y(n3723) );
  OAI21X1 U7139 ( .A(n12712), .B(n12821), .C(n3724), .Y(n7872) );
  NAND2X1 U7140 ( .A(ram[3435]), .B(n12821), .Y(n3724) );
  OAI21X1 U7141 ( .A(n12706), .B(n12821), .C(n3725), .Y(n7873) );
  NAND2X1 U7142 ( .A(ram[3436]), .B(n12821), .Y(n3725) );
  OAI21X1 U7143 ( .A(n12700), .B(n12821), .C(n3726), .Y(n7874) );
  NAND2X1 U7144 ( .A(ram[3437]), .B(n12821), .Y(n3726) );
  OAI21X1 U7145 ( .A(n12694), .B(n12821), .C(n3727), .Y(n7875) );
  NAND2X1 U7146 ( .A(ram[3438]), .B(n12821), .Y(n3727) );
  OAI21X1 U7147 ( .A(n12688), .B(n12821), .C(n3728), .Y(n7876) );
  NAND2X1 U7148 ( .A(ram[3439]), .B(n12821), .Y(n3728) );
  OAI21X1 U7150 ( .A(n12778), .B(n12820), .C(n3730), .Y(n7877) );
  NAND2X1 U7151 ( .A(ram[3440]), .B(n12820), .Y(n3730) );
  OAI21X1 U7152 ( .A(n12772), .B(n12820), .C(n3731), .Y(n7878) );
  NAND2X1 U7153 ( .A(ram[3441]), .B(n12820), .Y(n3731) );
  OAI21X1 U7154 ( .A(n12766), .B(n12820), .C(n3732), .Y(n7879) );
  NAND2X1 U7155 ( .A(ram[3442]), .B(n12820), .Y(n3732) );
  OAI21X1 U7156 ( .A(n12760), .B(n12820), .C(n3733), .Y(n7880) );
  NAND2X1 U7157 ( .A(ram[3443]), .B(n12820), .Y(n3733) );
  OAI21X1 U7158 ( .A(n12754), .B(n12820), .C(n3734), .Y(n7881) );
  NAND2X1 U7159 ( .A(ram[3444]), .B(n12820), .Y(n3734) );
  OAI21X1 U7160 ( .A(n12748), .B(n12820), .C(n3735), .Y(n7882) );
  NAND2X1 U7161 ( .A(ram[3445]), .B(n12820), .Y(n3735) );
  OAI21X1 U7162 ( .A(n12742), .B(n12820), .C(n3736), .Y(n7883) );
  NAND2X1 U7163 ( .A(ram[3446]), .B(n12820), .Y(n3736) );
  OAI21X1 U7164 ( .A(n12736), .B(n12820), .C(n3737), .Y(n7884) );
  NAND2X1 U7165 ( .A(ram[3447]), .B(n12820), .Y(n3737) );
  OAI21X1 U7166 ( .A(n12730), .B(n12820), .C(n3738), .Y(n7885) );
  NAND2X1 U7167 ( .A(ram[3448]), .B(n12820), .Y(n3738) );
  OAI21X1 U7168 ( .A(n12724), .B(n12820), .C(n3739), .Y(n7886) );
  NAND2X1 U7169 ( .A(ram[3449]), .B(n12820), .Y(n3739) );
  OAI21X1 U7170 ( .A(n12718), .B(n12820), .C(n3740), .Y(n7887) );
  NAND2X1 U7171 ( .A(ram[3450]), .B(n12820), .Y(n3740) );
  OAI21X1 U7172 ( .A(n12712), .B(n12820), .C(n3741), .Y(n7888) );
  NAND2X1 U7173 ( .A(ram[3451]), .B(n12820), .Y(n3741) );
  OAI21X1 U7174 ( .A(n12706), .B(n12820), .C(n3742), .Y(n7889) );
  NAND2X1 U7175 ( .A(ram[3452]), .B(n12820), .Y(n3742) );
  OAI21X1 U7176 ( .A(n12700), .B(n12820), .C(n3743), .Y(n7890) );
  NAND2X1 U7177 ( .A(ram[3453]), .B(n12820), .Y(n3743) );
  OAI21X1 U7178 ( .A(n12694), .B(n12820), .C(n3744), .Y(n7891) );
  NAND2X1 U7179 ( .A(ram[3454]), .B(n12820), .Y(n3744) );
  OAI21X1 U7180 ( .A(n12688), .B(n12820), .C(n3745), .Y(n7892) );
  NAND2X1 U7181 ( .A(ram[3455]), .B(n12820), .Y(n3745) );
  OAI21X1 U7183 ( .A(n12778), .B(n12819), .C(n3747), .Y(n7893) );
  NAND2X1 U7184 ( .A(ram[3456]), .B(n12819), .Y(n3747) );
  OAI21X1 U7185 ( .A(n12772), .B(n12819), .C(n3748), .Y(n7894) );
  NAND2X1 U7186 ( .A(ram[3457]), .B(n12819), .Y(n3748) );
  OAI21X1 U7187 ( .A(n12766), .B(n12819), .C(n3749), .Y(n7895) );
  NAND2X1 U7188 ( .A(ram[3458]), .B(n12819), .Y(n3749) );
  OAI21X1 U7189 ( .A(n12760), .B(n12819), .C(n3750), .Y(n7896) );
  NAND2X1 U7190 ( .A(ram[3459]), .B(n12819), .Y(n3750) );
  OAI21X1 U7191 ( .A(n12754), .B(n12819), .C(n3751), .Y(n7897) );
  NAND2X1 U7192 ( .A(ram[3460]), .B(n12819), .Y(n3751) );
  OAI21X1 U7193 ( .A(n12748), .B(n12819), .C(n3752), .Y(n7898) );
  NAND2X1 U7194 ( .A(ram[3461]), .B(n12819), .Y(n3752) );
  OAI21X1 U7195 ( .A(n12742), .B(n12819), .C(n3753), .Y(n7899) );
  NAND2X1 U7196 ( .A(ram[3462]), .B(n12819), .Y(n3753) );
  OAI21X1 U7197 ( .A(n12736), .B(n12819), .C(n3754), .Y(n7900) );
  NAND2X1 U7198 ( .A(ram[3463]), .B(n12819), .Y(n3754) );
  OAI21X1 U7199 ( .A(n12730), .B(n12819), .C(n3755), .Y(n7901) );
  NAND2X1 U7200 ( .A(ram[3464]), .B(n12819), .Y(n3755) );
  OAI21X1 U7201 ( .A(n12724), .B(n12819), .C(n3756), .Y(n7902) );
  NAND2X1 U7202 ( .A(ram[3465]), .B(n12819), .Y(n3756) );
  OAI21X1 U7203 ( .A(n12718), .B(n12819), .C(n3757), .Y(n7903) );
  NAND2X1 U7204 ( .A(ram[3466]), .B(n12819), .Y(n3757) );
  OAI21X1 U7205 ( .A(n12712), .B(n12819), .C(n3758), .Y(n7904) );
  NAND2X1 U7206 ( .A(ram[3467]), .B(n12819), .Y(n3758) );
  OAI21X1 U7207 ( .A(n12706), .B(n12819), .C(n3759), .Y(n7905) );
  NAND2X1 U7208 ( .A(ram[3468]), .B(n12819), .Y(n3759) );
  OAI21X1 U7209 ( .A(n12700), .B(n12819), .C(n3760), .Y(n7906) );
  NAND2X1 U7210 ( .A(ram[3469]), .B(n12819), .Y(n3760) );
  OAI21X1 U7211 ( .A(n12694), .B(n12819), .C(n3761), .Y(n7907) );
  NAND2X1 U7212 ( .A(ram[3470]), .B(n12819), .Y(n3761) );
  OAI21X1 U7213 ( .A(n12688), .B(n12819), .C(n3762), .Y(n7908) );
  NAND2X1 U7214 ( .A(ram[3471]), .B(n12819), .Y(n3762) );
  OAI21X1 U7216 ( .A(n12778), .B(n12818), .C(n3764), .Y(n7909) );
  NAND2X1 U7217 ( .A(ram[3472]), .B(n12818), .Y(n3764) );
  OAI21X1 U7218 ( .A(n12772), .B(n12818), .C(n3765), .Y(n7910) );
  NAND2X1 U7219 ( .A(ram[3473]), .B(n12818), .Y(n3765) );
  OAI21X1 U7220 ( .A(n12766), .B(n12818), .C(n3766), .Y(n7911) );
  NAND2X1 U7221 ( .A(ram[3474]), .B(n12818), .Y(n3766) );
  OAI21X1 U7222 ( .A(n12760), .B(n12818), .C(n3767), .Y(n7912) );
  NAND2X1 U7223 ( .A(ram[3475]), .B(n12818), .Y(n3767) );
  OAI21X1 U7224 ( .A(n12754), .B(n12818), .C(n3768), .Y(n7913) );
  NAND2X1 U7225 ( .A(ram[3476]), .B(n12818), .Y(n3768) );
  OAI21X1 U7226 ( .A(n12748), .B(n12818), .C(n3769), .Y(n7914) );
  NAND2X1 U7227 ( .A(ram[3477]), .B(n12818), .Y(n3769) );
  OAI21X1 U7228 ( .A(n12742), .B(n12818), .C(n3770), .Y(n7915) );
  NAND2X1 U7229 ( .A(ram[3478]), .B(n12818), .Y(n3770) );
  OAI21X1 U7230 ( .A(n12736), .B(n12818), .C(n3771), .Y(n7916) );
  NAND2X1 U7231 ( .A(ram[3479]), .B(n12818), .Y(n3771) );
  OAI21X1 U7232 ( .A(n12730), .B(n12818), .C(n3772), .Y(n7917) );
  NAND2X1 U7233 ( .A(ram[3480]), .B(n12818), .Y(n3772) );
  OAI21X1 U7234 ( .A(n12724), .B(n12818), .C(n3773), .Y(n7918) );
  NAND2X1 U7235 ( .A(ram[3481]), .B(n12818), .Y(n3773) );
  OAI21X1 U7236 ( .A(n12718), .B(n12818), .C(n3774), .Y(n7919) );
  NAND2X1 U7237 ( .A(ram[3482]), .B(n12818), .Y(n3774) );
  OAI21X1 U7238 ( .A(n12712), .B(n12818), .C(n3775), .Y(n7920) );
  NAND2X1 U7239 ( .A(ram[3483]), .B(n12818), .Y(n3775) );
  OAI21X1 U7240 ( .A(n12706), .B(n12818), .C(n3776), .Y(n7921) );
  NAND2X1 U7241 ( .A(ram[3484]), .B(n12818), .Y(n3776) );
  OAI21X1 U7242 ( .A(n12700), .B(n12818), .C(n3777), .Y(n7922) );
  NAND2X1 U7243 ( .A(ram[3485]), .B(n12818), .Y(n3777) );
  OAI21X1 U7244 ( .A(n12694), .B(n12818), .C(n3778), .Y(n7923) );
  NAND2X1 U7245 ( .A(ram[3486]), .B(n12818), .Y(n3778) );
  OAI21X1 U7246 ( .A(n12688), .B(n12818), .C(n3779), .Y(n7924) );
  NAND2X1 U7247 ( .A(ram[3487]), .B(n12818), .Y(n3779) );
  OAI21X1 U7249 ( .A(n12778), .B(n12817), .C(n3781), .Y(n7925) );
  NAND2X1 U7250 ( .A(ram[3488]), .B(n12817), .Y(n3781) );
  OAI21X1 U7251 ( .A(n12772), .B(n12817), .C(n3782), .Y(n7926) );
  NAND2X1 U7252 ( .A(ram[3489]), .B(n12817), .Y(n3782) );
  OAI21X1 U7253 ( .A(n12766), .B(n12817), .C(n3783), .Y(n7927) );
  NAND2X1 U7254 ( .A(ram[3490]), .B(n12817), .Y(n3783) );
  OAI21X1 U7255 ( .A(n12760), .B(n12817), .C(n3784), .Y(n7928) );
  NAND2X1 U7256 ( .A(ram[3491]), .B(n12817), .Y(n3784) );
  OAI21X1 U7257 ( .A(n12754), .B(n12817), .C(n3785), .Y(n7929) );
  NAND2X1 U7258 ( .A(ram[3492]), .B(n12817), .Y(n3785) );
  OAI21X1 U7259 ( .A(n12748), .B(n12817), .C(n3786), .Y(n7930) );
  NAND2X1 U7260 ( .A(ram[3493]), .B(n12817), .Y(n3786) );
  OAI21X1 U7261 ( .A(n12742), .B(n12817), .C(n3787), .Y(n7931) );
  NAND2X1 U7262 ( .A(ram[3494]), .B(n12817), .Y(n3787) );
  OAI21X1 U7263 ( .A(n12736), .B(n12817), .C(n3788), .Y(n7932) );
  NAND2X1 U7264 ( .A(ram[3495]), .B(n12817), .Y(n3788) );
  OAI21X1 U7265 ( .A(n12730), .B(n12817), .C(n3789), .Y(n7933) );
  NAND2X1 U7266 ( .A(ram[3496]), .B(n12817), .Y(n3789) );
  OAI21X1 U7267 ( .A(n12724), .B(n12817), .C(n3790), .Y(n7934) );
  NAND2X1 U7268 ( .A(ram[3497]), .B(n12817), .Y(n3790) );
  OAI21X1 U7269 ( .A(n12718), .B(n12817), .C(n3791), .Y(n7935) );
  NAND2X1 U7270 ( .A(ram[3498]), .B(n12817), .Y(n3791) );
  OAI21X1 U7271 ( .A(n12712), .B(n12817), .C(n3792), .Y(n7936) );
  NAND2X1 U7272 ( .A(ram[3499]), .B(n12817), .Y(n3792) );
  OAI21X1 U7273 ( .A(n12706), .B(n12817), .C(n3793), .Y(n7937) );
  NAND2X1 U7274 ( .A(ram[3500]), .B(n12817), .Y(n3793) );
  OAI21X1 U7275 ( .A(n12700), .B(n12817), .C(n3794), .Y(n7938) );
  NAND2X1 U7276 ( .A(ram[3501]), .B(n12817), .Y(n3794) );
  OAI21X1 U7277 ( .A(n12694), .B(n12817), .C(n3795), .Y(n7939) );
  NAND2X1 U7278 ( .A(ram[3502]), .B(n12817), .Y(n3795) );
  OAI21X1 U7279 ( .A(n12688), .B(n12817), .C(n3796), .Y(n7940) );
  NAND2X1 U7280 ( .A(ram[3503]), .B(n12817), .Y(n3796) );
  OAI21X1 U7282 ( .A(n12778), .B(n12816), .C(n3798), .Y(n7941) );
  NAND2X1 U7283 ( .A(ram[3504]), .B(n12816), .Y(n3798) );
  OAI21X1 U7284 ( .A(n12772), .B(n12816), .C(n3799), .Y(n7942) );
  NAND2X1 U7285 ( .A(ram[3505]), .B(n12816), .Y(n3799) );
  OAI21X1 U7286 ( .A(n12766), .B(n12816), .C(n3800), .Y(n7943) );
  NAND2X1 U7287 ( .A(ram[3506]), .B(n12816), .Y(n3800) );
  OAI21X1 U7288 ( .A(n12760), .B(n12816), .C(n3801), .Y(n7944) );
  NAND2X1 U7289 ( .A(ram[3507]), .B(n12816), .Y(n3801) );
  OAI21X1 U7290 ( .A(n12754), .B(n12816), .C(n3802), .Y(n7945) );
  NAND2X1 U7291 ( .A(ram[3508]), .B(n12816), .Y(n3802) );
  OAI21X1 U7292 ( .A(n12748), .B(n12816), .C(n3803), .Y(n7946) );
  NAND2X1 U7293 ( .A(ram[3509]), .B(n12816), .Y(n3803) );
  OAI21X1 U7294 ( .A(n12742), .B(n12816), .C(n3804), .Y(n7947) );
  NAND2X1 U7295 ( .A(ram[3510]), .B(n12816), .Y(n3804) );
  OAI21X1 U7296 ( .A(n12736), .B(n12816), .C(n3805), .Y(n7948) );
  NAND2X1 U7297 ( .A(ram[3511]), .B(n12816), .Y(n3805) );
  OAI21X1 U7298 ( .A(n12730), .B(n12816), .C(n3806), .Y(n7949) );
  NAND2X1 U7299 ( .A(ram[3512]), .B(n12816), .Y(n3806) );
  OAI21X1 U7300 ( .A(n12724), .B(n12816), .C(n3807), .Y(n7950) );
  NAND2X1 U7301 ( .A(ram[3513]), .B(n12816), .Y(n3807) );
  OAI21X1 U7302 ( .A(n12718), .B(n12816), .C(n3808), .Y(n7951) );
  NAND2X1 U7303 ( .A(ram[3514]), .B(n12816), .Y(n3808) );
  OAI21X1 U7304 ( .A(n12712), .B(n12816), .C(n3809), .Y(n7952) );
  NAND2X1 U7305 ( .A(ram[3515]), .B(n12816), .Y(n3809) );
  OAI21X1 U7306 ( .A(n12706), .B(n12816), .C(n3810), .Y(n7953) );
  NAND2X1 U7307 ( .A(ram[3516]), .B(n12816), .Y(n3810) );
  OAI21X1 U7308 ( .A(n12700), .B(n12816), .C(n3811), .Y(n7954) );
  NAND2X1 U7309 ( .A(ram[3517]), .B(n12816), .Y(n3811) );
  OAI21X1 U7310 ( .A(n12694), .B(n12816), .C(n3812), .Y(n7955) );
  NAND2X1 U7311 ( .A(ram[3518]), .B(n12816), .Y(n3812) );
  OAI21X1 U7312 ( .A(n12688), .B(n12816), .C(n3813), .Y(n7956) );
  NAND2X1 U7313 ( .A(ram[3519]), .B(n12816), .Y(n3813) );
  OAI21X1 U7315 ( .A(n12778), .B(n12815), .C(n3815), .Y(n7957) );
  NAND2X1 U7316 ( .A(ram[3520]), .B(n12815), .Y(n3815) );
  OAI21X1 U7317 ( .A(n12772), .B(n12815), .C(n3816), .Y(n7958) );
  NAND2X1 U7318 ( .A(ram[3521]), .B(n12815), .Y(n3816) );
  OAI21X1 U7319 ( .A(n12766), .B(n12815), .C(n3817), .Y(n7959) );
  NAND2X1 U7320 ( .A(ram[3522]), .B(n12815), .Y(n3817) );
  OAI21X1 U7321 ( .A(n12760), .B(n12815), .C(n3818), .Y(n7960) );
  NAND2X1 U7322 ( .A(ram[3523]), .B(n12815), .Y(n3818) );
  OAI21X1 U7323 ( .A(n12754), .B(n12815), .C(n3819), .Y(n7961) );
  NAND2X1 U7324 ( .A(ram[3524]), .B(n12815), .Y(n3819) );
  OAI21X1 U7325 ( .A(n12748), .B(n12815), .C(n3820), .Y(n7962) );
  NAND2X1 U7326 ( .A(ram[3525]), .B(n12815), .Y(n3820) );
  OAI21X1 U7327 ( .A(n12742), .B(n12815), .C(n3821), .Y(n7963) );
  NAND2X1 U7328 ( .A(ram[3526]), .B(n12815), .Y(n3821) );
  OAI21X1 U7329 ( .A(n12736), .B(n12815), .C(n3822), .Y(n7964) );
  NAND2X1 U7330 ( .A(ram[3527]), .B(n12815), .Y(n3822) );
  OAI21X1 U7331 ( .A(n12730), .B(n12815), .C(n3823), .Y(n7965) );
  NAND2X1 U7332 ( .A(ram[3528]), .B(n12815), .Y(n3823) );
  OAI21X1 U7333 ( .A(n12724), .B(n12815), .C(n3824), .Y(n7966) );
  NAND2X1 U7334 ( .A(ram[3529]), .B(n12815), .Y(n3824) );
  OAI21X1 U7335 ( .A(n12718), .B(n12815), .C(n3825), .Y(n7967) );
  NAND2X1 U7336 ( .A(ram[3530]), .B(n12815), .Y(n3825) );
  OAI21X1 U7337 ( .A(n12712), .B(n12815), .C(n3826), .Y(n7968) );
  NAND2X1 U7338 ( .A(ram[3531]), .B(n12815), .Y(n3826) );
  OAI21X1 U7339 ( .A(n12706), .B(n12815), .C(n3827), .Y(n7969) );
  NAND2X1 U7340 ( .A(ram[3532]), .B(n12815), .Y(n3827) );
  OAI21X1 U7341 ( .A(n12700), .B(n12815), .C(n3828), .Y(n7970) );
  NAND2X1 U7342 ( .A(ram[3533]), .B(n12815), .Y(n3828) );
  OAI21X1 U7343 ( .A(n12694), .B(n12815), .C(n3829), .Y(n7971) );
  NAND2X1 U7344 ( .A(ram[3534]), .B(n12815), .Y(n3829) );
  OAI21X1 U7345 ( .A(n12688), .B(n12815), .C(n3830), .Y(n7972) );
  NAND2X1 U7346 ( .A(ram[3535]), .B(n12815), .Y(n3830) );
  OAI21X1 U7348 ( .A(n12779), .B(n12814), .C(n3832), .Y(n7973) );
  NAND2X1 U7349 ( .A(ram[3536]), .B(n12814), .Y(n3832) );
  OAI21X1 U7350 ( .A(n12773), .B(n12814), .C(n3833), .Y(n7974) );
  NAND2X1 U7351 ( .A(ram[3537]), .B(n12814), .Y(n3833) );
  OAI21X1 U7352 ( .A(n12767), .B(n12814), .C(n3834), .Y(n7975) );
  NAND2X1 U7353 ( .A(ram[3538]), .B(n12814), .Y(n3834) );
  OAI21X1 U7354 ( .A(n12761), .B(n12814), .C(n3835), .Y(n7976) );
  NAND2X1 U7355 ( .A(ram[3539]), .B(n12814), .Y(n3835) );
  OAI21X1 U7356 ( .A(n12755), .B(n12814), .C(n3836), .Y(n7977) );
  NAND2X1 U7357 ( .A(ram[3540]), .B(n12814), .Y(n3836) );
  OAI21X1 U7358 ( .A(n12749), .B(n12814), .C(n3837), .Y(n7978) );
  NAND2X1 U7359 ( .A(ram[3541]), .B(n12814), .Y(n3837) );
  OAI21X1 U7360 ( .A(n12743), .B(n12814), .C(n3838), .Y(n7979) );
  NAND2X1 U7361 ( .A(ram[3542]), .B(n12814), .Y(n3838) );
  OAI21X1 U7362 ( .A(n12737), .B(n12814), .C(n3839), .Y(n7980) );
  NAND2X1 U7363 ( .A(ram[3543]), .B(n12814), .Y(n3839) );
  OAI21X1 U7364 ( .A(n12731), .B(n12814), .C(n3840), .Y(n7981) );
  NAND2X1 U7365 ( .A(ram[3544]), .B(n12814), .Y(n3840) );
  OAI21X1 U7366 ( .A(n12725), .B(n12814), .C(n3841), .Y(n7982) );
  NAND2X1 U7367 ( .A(ram[3545]), .B(n12814), .Y(n3841) );
  OAI21X1 U7368 ( .A(n12719), .B(n12814), .C(n3842), .Y(n7983) );
  NAND2X1 U7369 ( .A(ram[3546]), .B(n12814), .Y(n3842) );
  OAI21X1 U7370 ( .A(n12713), .B(n12814), .C(n3843), .Y(n7984) );
  NAND2X1 U7371 ( .A(ram[3547]), .B(n12814), .Y(n3843) );
  OAI21X1 U7372 ( .A(n12707), .B(n12814), .C(n3844), .Y(n7985) );
  NAND2X1 U7373 ( .A(ram[3548]), .B(n12814), .Y(n3844) );
  OAI21X1 U7374 ( .A(n12701), .B(n12814), .C(n3845), .Y(n7986) );
  NAND2X1 U7375 ( .A(ram[3549]), .B(n12814), .Y(n3845) );
  OAI21X1 U7376 ( .A(n12695), .B(n12814), .C(n3846), .Y(n7987) );
  NAND2X1 U7377 ( .A(ram[3550]), .B(n12814), .Y(n3846) );
  OAI21X1 U7378 ( .A(n12689), .B(n12814), .C(n3847), .Y(n7988) );
  NAND2X1 U7379 ( .A(ram[3551]), .B(n12814), .Y(n3847) );
  OAI21X1 U7381 ( .A(n12779), .B(n12813), .C(n3849), .Y(n7989) );
  NAND2X1 U7382 ( .A(ram[3552]), .B(n12813), .Y(n3849) );
  OAI21X1 U7383 ( .A(n12773), .B(n12813), .C(n3850), .Y(n7990) );
  NAND2X1 U7384 ( .A(ram[3553]), .B(n12813), .Y(n3850) );
  OAI21X1 U7385 ( .A(n12767), .B(n12813), .C(n3851), .Y(n7991) );
  NAND2X1 U7386 ( .A(ram[3554]), .B(n12813), .Y(n3851) );
  OAI21X1 U7387 ( .A(n12761), .B(n12813), .C(n3852), .Y(n7992) );
  NAND2X1 U7388 ( .A(ram[3555]), .B(n12813), .Y(n3852) );
  OAI21X1 U7389 ( .A(n12755), .B(n12813), .C(n3853), .Y(n7993) );
  NAND2X1 U7390 ( .A(ram[3556]), .B(n12813), .Y(n3853) );
  OAI21X1 U7391 ( .A(n12749), .B(n12813), .C(n3854), .Y(n7994) );
  NAND2X1 U7392 ( .A(ram[3557]), .B(n12813), .Y(n3854) );
  OAI21X1 U7393 ( .A(n12743), .B(n12813), .C(n3855), .Y(n7995) );
  NAND2X1 U7394 ( .A(ram[3558]), .B(n12813), .Y(n3855) );
  OAI21X1 U7395 ( .A(n12737), .B(n12813), .C(n3856), .Y(n7996) );
  NAND2X1 U7396 ( .A(ram[3559]), .B(n12813), .Y(n3856) );
  OAI21X1 U7397 ( .A(n12731), .B(n12813), .C(n3857), .Y(n7997) );
  NAND2X1 U7398 ( .A(ram[3560]), .B(n12813), .Y(n3857) );
  OAI21X1 U7399 ( .A(n12725), .B(n12813), .C(n3858), .Y(n7998) );
  NAND2X1 U7400 ( .A(ram[3561]), .B(n12813), .Y(n3858) );
  OAI21X1 U7401 ( .A(n12719), .B(n12813), .C(n3859), .Y(n7999) );
  NAND2X1 U7402 ( .A(ram[3562]), .B(n12813), .Y(n3859) );
  OAI21X1 U7403 ( .A(n12713), .B(n12813), .C(n3860), .Y(n8000) );
  NAND2X1 U7404 ( .A(ram[3563]), .B(n12813), .Y(n3860) );
  OAI21X1 U7405 ( .A(n12707), .B(n12813), .C(n3861), .Y(n8001) );
  NAND2X1 U7406 ( .A(ram[3564]), .B(n12813), .Y(n3861) );
  OAI21X1 U7407 ( .A(n12701), .B(n12813), .C(n3862), .Y(n8002) );
  NAND2X1 U7408 ( .A(ram[3565]), .B(n12813), .Y(n3862) );
  OAI21X1 U7409 ( .A(n12695), .B(n12813), .C(n3863), .Y(n8003) );
  NAND2X1 U7410 ( .A(ram[3566]), .B(n12813), .Y(n3863) );
  OAI21X1 U7411 ( .A(n12689), .B(n12813), .C(n3864), .Y(n8004) );
  NAND2X1 U7412 ( .A(ram[3567]), .B(n12813), .Y(n3864) );
  OAI21X1 U7414 ( .A(n12779), .B(n12812), .C(n3866), .Y(n8005) );
  NAND2X1 U7415 ( .A(ram[3568]), .B(n12812), .Y(n3866) );
  OAI21X1 U7416 ( .A(n12773), .B(n12812), .C(n3867), .Y(n8006) );
  NAND2X1 U7417 ( .A(ram[3569]), .B(n12812), .Y(n3867) );
  OAI21X1 U7418 ( .A(n12767), .B(n12812), .C(n3868), .Y(n8007) );
  NAND2X1 U7419 ( .A(ram[3570]), .B(n12812), .Y(n3868) );
  OAI21X1 U7420 ( .A(n12761), .B(n12812), .C(n3869), .Y(n8008) );
  NAND2X1 U7421 ( .A(ram[3571]), .B(n12812), .Y(n3869) );
  OAI21X1 U7422 ( .A(n12755), .B(n12812), .C(n3870), .Y(n8009) );
  NAND2X1 U7423 ( .A(ram[3572]), .B(n12812), .Y(n3870) );
  OAI21X1 U7424 ( .A(n12749), .B(n12812), .C(n3871), .Y(n8010) );
  NAND2X1 U7425 ( .A(ram[3573]), .B(n12812), .Y(n3871) );
  OAI21X1 U7426 ( .A(n12743), .B(n12812), .C(n3872), .Y(n8011) );
  NAND2X1 U7427 ( .A(ram[3574]), .B(n12812), .Y(n3872) );
  OAI21X1 U7428 ( .A(n12737), .B(n12812), .C(n3873), .Y(n8012) );
  NAND2X1 U7429 ( .A(ram[3575]), .B(n12812), .Y(n3873) );
  OAI21X1 U7430 ( .A(n12731), .B(n12812), .C(n3874), .Y(n8013) );
  NAND2X1 U7431 ( .A(ram[3576]), .B(n12812), .Y(n3874) );
  OAI21X1 U7432 ( .A(n12725), .B(n12812), .C(n3875), .Y(n8014) );
  NAND2X1 U7433 ( .A(ram[3577]), .B(n12812), .Y(n3875) );
  OAI21X1 U7434 ( .A(n12719), .B(n12812), .C(n3876), .Y(n8015) );
  NAND2X1 U7435 ( .A(ram[3578]), .B(n12812), .Y(n3876) );
  OAI21X1 U7436 ( .A(n12713), .B(n12812), .C(n3877), .Y(n8016) );
  NAND2X1 U7437 ( .A(ram[3579]), .B(n12812), .Y(n3877) );
  OAI21X1 U7438 ( .A(n12707), .B(n12812), .C(n3878), .Y(n8017) );
  NAND2X1 U7439 ( .A(ram[3580]), .B(n12812), .Y(n3878) );
  OAI21X1 U7440 ( .A(n12701), .B(n12812), .C(n3879), .Y(n8018) );
  NAND2X1 U7441 ( .A(ram[3581]), .B(n12812), .Y(n3879) );
  OAI21X1 U7442 ( .A(n12695), .B(n12812), .C(n3880), .Y(n8019) );
  NAND2X1 U7443 ( .A(ram[3582]), .B(n12812), .Y(n3880) );
  OAI21X1 U7444 ( .A(n12689), .B(n12812), .C(n3881), .Y(n8020) );
  NAND2X1 U7445 ( .A(ram[3583]), .B(n12812), .Y(n3881) );
  NAND3X1 U7447 ( .A(n601), .B(mem_write_en), .C(n3609), .Y(n3882) );
  NOR2X1 U7448 ( .A(n13038), .B(mem_access_addr[5]), .Y(n601) );
  OAI21X1 U7449 ( .A(n12779), .B(n12811), .C(n3884), .Y(n8021) );
  NAND2X1 U7450 ( .A(ram[3584]), .B(n12811), .Y(n3884) );
  OAI21X1 U7451 ( .A(n12773), .B(n12811), .C(n3885), .Y(n8022) );
  NAND2X1 U7452 ( .A(ram[3585]), .B(n12811), .Y(n3885) );
  OAI21X1 U7453 ( .A(n12767), .B(n12811), .C(n3886), .Y(n8023) );
  NAND2X1 U7454 ( .A(ram[3586]), .B(n12811), .Y(n3886) );
  OAI21X1 U7455 ( .A(n12761), .B(n12811), .C(n3887), .Y(n8024) );
  NAND2X1 U7456 ( .A(ram[3587]), .B(n12811), .Y(n3887) );
  OAI21X1 U7457 ( .A(n12755), .B(n12811), .C(n3888), .Y(n8025) );
  NAND2X1 U7458 ( .A(ram[3588]), .B(n12811), .Y(n3888) );
  OAI21X1 U7459 ( .A(n12749), .B(n12811), .C(n3889), .Y(n8026) );
  NAND2X1 U7460 ( .A(ram[3589]), .B(n12811), .Y(n3889) );
  OAI21X1 U7461 ( .A(n12743), .B(n12811), .C(n3890), .Y(n8027) );
  NAND2X1 U7462 ( .A(ram[3590]), .B(n12811), .Y(n3890) );
  OAI21X1 U7463 ( .A(n12737), .B(n12811), .C(n3891), .Y(n8028) );
  NAND2X1 U7464 ( .A(ram[3591]), .B(n12811), .Y(n3891) );
  OAI21X1 U7465 ( .A(n12731), .B(n12811), .C(n3892), .Y(n8029) );
  NAND2X1 U7466 ( .A(ram[3592]), .B(n12811), .Y(n3892) );
  OAI21X1 U7467 ( .A(n12725), .B(n12811), .C(n3893), .Y(n8030) );
  NAND2X1 U7468 ( .A(ram[3593]), .B(n12811), .Y(n3893) );
  OAI21X1 U7469 ( .A(n12719), .B(n12811), .C(n3894), .Y(n8031) );
  NAND2X1 U7470 ( .A(ram[3594]), .B(n12811), .Y(n3894) );
  OAI21X1 U7471 ( .A(n12713), .B(n12811), .C(n3895), .Y(n8032) );
  NAND2X1 U7472 ( .A(ram[3595]), .B(n12811), .Y(n3895) );
  OAI21X1 U7473 ( .A(n12707), .B(n12811), .C(n3896), .Y(n8033) );
  NAND2X1 U7474 ( .A(ram[3596]), .B(n12811), .Y(n3896) );
  OAI21X1 U7475 ( .A(n12701), .B(n12811), .C(n3897), .Y(n8034) );
  NAND2X1 U7476 ( .A(ram[3597]), .B(n12811), .Y(n3897) );
  OAI21X1 U7477 ( .A(n12695), .B(n12811), .C(n3898), .Y(n8035) );
  NAND2X1 U7478 ( .A(ram[3598]), .B(n12811), .Y(n3898) );
  OAI21X1 U7479 ( .A(n12689), .B(n12811), .C(n3899), .Y(n8036) );
  NAND2X1 U7480 ( .A(ram[3599]), .B(n12811), .Y(n3899) );
  OAI21X1 U7482 ( .A(n12779), .B(n12810), .C(n3901), .Y(n8037) );
  NAND2X1 U7483 ( .A(ram[3600]), .B(n12810), .Y(n3901) );
  OAI21X1 U7484 ( .A(n12773), .B(n12810), .C(n3902), .Y(n8038) );
  NAND2X1 U7485 ( .A(ram[3601]), .B(n12810), .Y(n3902) );
  OAI21X1 U7486 ( .A(n12767), .B(n12810), .C(n3903), .Y(n8039) );
  NAND2X1 U7487 ( .A(ram[3602]), .B(n12810), .Y(n3903) );
  OAI21X1 U7488 ( .A(n12761), .B(n12810), .C(n3904), .Y(n8040) );
  NAND2X1 U7489 ( .A(ram[3603]), .B(n12810), .Y(n3904) );
  OAI21X1 U7490 ( .A(n12755), .B(n12810), .C(n3905), .Y(n8041) );
  NAND2X1 U7491 ( .A(ram[3604]), .B(n12810), .Y(n3905) );
  OAI21X1 U7492 ( .A(n12749), .B(n12810), .C(n3906), .Y(n8042) );
  NAND2X1 U7493 ( .A(ram[3605]), .B(n12810), .Y(n3906) );
  OAI21X1 U7494 ( .A(n12743), .B(n12810), .C(n3907), .Y(n8043) );
  NAND2X1 U7495 ( .A(ram[3606]), .B(n12810), .Y(n3907) );
  OAI21X1 U7496 ( .A(n12737), .B(n12810), .C(n3908), .Y(n8044) );
  NAND2X1 U7497 ( .A(ram[3607]), .B(n12810), .Y(n3908) );
  OAI21X1 U7498 ( .A(n12731), .B(n12810), .C(n3909), .Y(n8045) );
  NAND2X1 U7499 ( .A(ram[3608]), .B(n12810), .Y(n3909) );
  OAI21X1 U7500 ( .A(n12725), .B(n12810), .C(n3910), .Y(n8046) );
  NAND2X1 U7501 ( .A(ram[3609]), .B(n12810), .Y(n3910) );
  OAI21X1 U7502 ( .A(n12719), .B(n12810), .C(n3911), .Y(n8047) );
  NAND2X1 U7503 ( .A(ram[3610]), .B(n12810), .Y(n3911) );
  OAI21X1 U7504 ( .A(n12713), .B(n12810), .C(n3912), .Y(n8048) );
  NAND2X1 U7505 ( .A(ram[3611]), .B(n12810), .Y(n3912) );
  OAI21X1 U7506 ( .A(n12707), .B(n12810), .C(n3913), .Y(n8049) );
  NAND2X1 U7507 ( .A(ram[3612]), .B(n12810), .Y(n3913) );
  OAI21X1 U7508 ( .A(n12701), .B(n12810), .C(n3914), .Y(n8050) );
  NAND2X1 U7509 ( .A(ram[3613]), .B(n12810), .Y(n3914) );
  OAI21X1 U7510 ( .A(n12695), .B(n12810), .C(n3915), .Y(n8051) );
  NAND2X1 U7511 ( .A(ram[3614]), .B(n12810), .Y(n3915) );
  OAI21X1 U7512 ( .A(n12689), .B(n12810), .C(n3916), .Y(n8052) );
  NAND2X1 U7513 ( .A(ram[3615]), .B(n12810), .Y(n3916) );
  OAI21X1 U7515 ( .A(n12779), .B(n12809), .C(n3918), .Y(n8053) );
  NAND2X1 U7516 ( .A(ram[3616]), .B(n12809), .Y(n3918) );
  OAI21X1 U7517 ( .A(n12773), .B(n12809), .C(n3919), .Y(n8054) );
  NAND2X1 U7518 ( .A(ram[3617]), .B(n12809), .Y(n3919) );
  OAI21X1 U7519 ( .A(n12767), .B(n12809), .C(n3920), .Y(n8055) );
  NAND2X1 U7520 ( .A(ram[3618]), .B(n12809), .Y(n3920) );
  OAI21X1 U7521 ( .A(n12761), .B(n12809), .C(n3921), .Y(n8056) );
  NAND2X1 U7522 ( .A(ram[3619]), .B(n12809), .Y(n3921) );
  OAI21X1 U7523 ( .A(n12755), .B(n12809), .C(n3922), .Y(n8057) );
  NAND2X1 U7524 ( .A(ram[3620]), .B(n12809), .Y(n3922) );
  OAI21X1 U7525 ( .A(n12749), .B(n12809), .C(n3923), .Y(n8058) );
  NAND2X1 U7526 ( .A(ram[3621]), .B(n12809), .Y(n3923) );
  OAI21X1 U7527 ( .A(n12743), .B(n12809), .C(n3924), .Y(n8059) );
  NAND2X1 U7528 ( .A(ram[3622]), .B(n12809), .Y(n3924) );
  OAI21X1 U7529 ( .A(n12737), .B(n12809), .C(n3925), .Y(n8060) );
  NAND2X1 U7530 ( .A(ram[3623]), .B(n12809), .Y(n3925) );
  OAI21X1 U7531 ( .A(n12731), .B(n12809), .C(n3926), .Y(n8061) );
  NAND2X1 U7532 ( .A(ram[3624]), .B(n12809), .Y(n3926) );
  OAI21X1 U7533 ( .A(n12725), .B(n12809), .C(n3927), .Y(n8062) );
  NAND2X1 U7534 ( .A(ram[3625]), .B(n12809), .Y(n3927) );
  OAI21X1 U7535 ( .A(n12719), .B(n12809), .C(n3928), .Y(n8063) );
  NAND2X1 U7536 ( .A(ram[3626]), .B(n12809), .Y(n3928) );
  OAI21X1 U7537 ( .A(n12713), .B(n12809), .C(n3929), .Y(n8064) );
  NAND2X1 U7538 ( .A(ram[3627]), .B(n12809), .Y(n3929) );
  OAI21X1 U7539 ( .A(n12707), .B(n12809), .C(n3930), .Y(n8065) );
  NAND2X1 U7540 ( .A(ram[3628]), .B(n12809), .Y(n3930) );
  OAI21X1 U7541 ( .A(n12701), .B(n12809), .C(n3931), .Y(n8066) );
  NAND2X1 U7542 ( .A(ram[3629]), .B(n12809), .Y(n3931) );
  OAI21X1 U7543 ( .A(n12695), .B(n12809), .C(n3932), .Y(n8067) );
  NAND2X1 U7544 ( .A(ram[3630]), .B(n12809), .Y(n3932) );
  OAI21X1 U7545 ( .A(n12689), .B(n12809), .C(n3933), .Y(n8068) );
  NAND2X1 U7546 ( .A(ram[3631]), .B(n12809), .Y(n3933) );
  OAI21X1 U7548 ( .A(n12779), .B(n12808), .C(n3935), .Y(n8069) );
  NAND2X1 U7549 ( .A(ram[3632]), .B(n12808), .Y(n3935) );
  OAI21X1 U7550 ( .A(n12773), .B(n12808), .C(n3936), .Y(n8070) );
  NAND2X1 U7551 ( .A(ram[3633]), .B(n12808), .Y(n3936) );
  OAI21X1 U7552 ( .A(n12767), .B(n12808), .C(n3937), .Y(n8071) );
  NAND2X1 U7553 ( .A(ram[3634]), .B(n12808), .Y(n3937) );
  OAI21X1 U7554 ( .A(n12761), .B(n12808), .C(n3938), .Y(n8072) );
  NAND2X1 U7555 ( .A(ram[3635]), .B(n12808), .Y(n3938) );
  OAI21X1 U7556 ( .A(n12755), .B(n12808), .C(n3939), .Y(n8073) );
  NAND2X1 U7557 ( .A(ram[3636]), .B(n12808), .Y(n3939) );
  OAI21X1 U7558 ( .A(n12749), .B(n12808), .C(n3940), .Y(n8074) );
  NAND2X1 U7559 ( .A(ram[3637]), .B(n12808), .Y(n3940) );
  OAI21X1 U7560 ( .A(n12743), .B(n12808), .C(n3941), .Y(n8075) );
  NAND2X1 U7561 ( .A(ram[3638]), .B(n12808), .Y(n3941) );
  OAI21X1 U7562 ( .A(n12737), .B(n12808), .C(n3942), .Y(n8076) );
  NAND2X1 U7563 ( .A(ram[3639]), .B(n12808), .Y(n3942) );
  OAI21X1 U7564 ( .A(n12731), .B(n12808), .C(n3943), .Y(n8077) );
  NAND2X1 U7565 ( .A(ram[3640]), .B(n12808), .Y(n3943) );
  OAI21X1 U7566 ( .A(n12725), .B(n12808), .C(n3944), .Y(n8078) );
  NAND2X1 U7567 ( .A(ram[3641]), .B(n12808), .Y(n3944) );
  OAI21X1 U7568 ( .A(n12719), .B(n12808), .C(n3945), .Y(n8079) );
  NAND2X1 U7569 ( .A(ram[3642]), .B(n12808), .Y(n3945) );
  OAI21X1 U7570 ( .A(n12713), .B(n12808), .C(n3946), .Y(n8080) );
  NAND2X1 U7571 ( .A(ram[3643]), .B(n12808), .Y(n3946) );
  OAI21X1 U7572 ( .A(n12707), .B(n12808), .C(n3947), .Y(n8081) );
  NAND2X1 U7573 ( .A(ram[3644]), .B(n12808), .Y(n3947) );
  OAI21X1 U7574 ( .A(n12701), .B(n12808), .C(n3948), .Y(n8082) );
  NAND2X1 U7575 ( .A(ram[3645]), .B(n12808), .Y(n3948) );
  OAI21X1 U7576 ( .A(n12695), .B(n12808), .C(n3949), .Y(n8083) );
  NAND2X1 U7577 ( .A(ram[3646]), .B(n12808), .Y(n3949) );
  OAI21X1 U7578 ( .A(n12689), .B(n12808), .C(n3950), .Y(n8084) );
  NAND2X1 U7579 ( .A(ram[3647]), .B(n12808), .Y(n3950) );
  OAI21X1 U7581 ( .A(n12779), .B(n12807), .C(n3952), .Y(n8085) );
  NAND2X1 U7582 ( .A(ram[3648]), .B(n12807), .Y(n3952) );
  OAI21X1 U7583 ( .A(n12773), .B(n12807), .C(n3953), .Y(n8086) );
  NAND2X1 U7584 ( .A(ram[3649]), .B(n12807), .Y(n3953) );
  OAI21X1 U7585 ( .A(n12767), .B(n12807), .C(n3954), .Y(n8087) );
  NAND2X1 U7586 ( .A(ram[3650]), .B(n12807), .Y(n3954) );
  OAI21X1 U7587 ( .A(n12761), .B(n12807), .C(n3955), .Y(n8088) );
  NAND2X1 U7588 ( .A(ram[3651]), .B(n12807), .Y(n3955) );
  OAI21X1 U7589 ( .A(n12755), .B(n12807), .C(n3956), .Y(n8089) );
  NAND2X1 U7590 ( .A(ram[3652]), .B(n12807), .Y(n3956) );
  OAI21X1 U7591 ( .A(n12749), .B(n12807), .C(n3957), .Y(n8090) );
  NAND2X1 U7592 ( .A(ram[3653]), .B(n12807), .Y(n3957) );
  OAI21X1 U7593 ( .A(n12743), .B(n12807), .C(n3958), .Y(n8091) );
  NAND2X1 U7594 ( .A(ram[3654]), .B(n12807), .Y(n3958) );
  OAI21X1 U7595 ( .A(n12737), .B(n12807), .C(n3959), .Y(n8092) );
  NAND2X1 U7596 ( .A(ram[3655]), .B(n12807), .Y(n3959) );
  OAI21X1 U7597 ( .A(n12731), .B(n12807), .C(n3960), .Y(n8093) );
  NAND2X1 U7598 ( .A(ram[3656]), .B(n12807), .Y(n3960) );
  OAI21X1 U7599 ( .A(n12725), .B(n12807), .C(n3961), .Y(n8094) );
  NAND2X1 U7600 ( .A(ram[3657]), .B(n12807), .Y(n3961) );
  OAI21X1 U7601 ( .A(n12719), .B(n12807), .C(n3962), .Y(n8095) );
  NAND2X1 U7602 ( .A(ram[3658]), .B(n12807), .Y(n3962) );
  OAI21X1 U7603 ( .A(n12713), .B(n12807), .C(n3963), .Y(n8096) );
  NAND2X1 U7604 ( .A(ram[3659]), .B(n12807), .Y(n3963) );
  OAI21X1 U7605 ( .A(n12707), .B(n12807), .C(n3964), .Y(n8097) );
  NAND2X1 U7606 ( .A(ram[3660]), .B(n12807), .Y(n3964) );
  OAI21X1 U7607 ( .A(n12701), .B(n12807), .C(n3965), .Y(n8098) );
  NAND2X1 U7608 ( .A(ram[3661]), .B(n12807), .Y(n3965) );
  OAI21X1 U7609 ( .A(n12695), .B(n12807), .C(n3966), .Y(n8099) );
  NAND2X1 U7610 ( .A(ram[3662]), .B(n12807), .Y(n3966) );
  OAI21X1 U7611 ( .A(n12689), .B(n12807), .C(n3967), .Y(n8100) );
  NAND2X1 U7612 ( .A(ram[3663]), .B(n12807), .Y(n3967) );
  OAI21X1 U7614 ( .A(n12779), .B(n12806), .C(n3969), .Y(n8101) );
  NAND2X1 U7615 ( .A(ram[3664]), .B(n12806), .Y(n3969) );
  OAI21X1 U7616 ( .A(n12773), .B(n12806), .C(n3970), .Y(n8102) );
  NAND2X1 U7617 ( .A(ram[3665]), .B(n12806), .Y(n3970) );
  OAI21X1 U7618 ( .A(n12767), .B(n12806), .C(n3971), .Y(n8103) );
  NAND2X1 U7619 ( .A(ram[3666]), .B(n12806), .Y(n3971) );
  OAI21X1 U7620 ( .A(n12761), .B(n12806), .C(n3972), .Y(n8104) );
  NAND2X1 U7621 ( .A(ram[3667]), .B(n12806), .Y(n3972) );
  OAI21X1 U7622 ( .A(n12755), .B(n12806), .C(n3973), .Y(n8105) );
  NAND2X1 U7623 ( .A(ram[3668]), .B(n12806), .Y(n3973) );
  OAI21X1 U7624 ( .A(n12749), .B(n12806), .C(n3974), .Y(n8106) );
  NAND2X1 U7625 ( .A(ram[3669]), .B(n12806), .Y(n3974) );
  OAI21X1 U7626 ( .A(n12743), .B(n12806), .C(n3975), .Y(n8107) );
  NAND2X1 U7627 ( .A(ram[3670]), .B(n12806), .Y(n3975) );
  OAI21X1 U7628 ( .A(n12737), .B(n12806), .C(n3976), .Y(n8108) );
  NAND2X1 U7629 ( .A(ram[3671]), .B(n12806), .Y(n3976) );
  OAI21X1 U7630 ( .A(n12731), .B(n12806), .C(n3977), .Y(n8109) );
  NAND2X1 U7631 ( .A(ram[3672]), .B(n12806), .Y(n3977) );
  OAI21X1 U7632 ( .A(n12725), .B(n12806), .C(n3978), .Y(n8110) );
  NAND2X1 U7633 ( .A(ram[3673]), .B(n12806), .Y(n3978) );
  OAI21X1 U7634 ( .A(n12719), .B(n12806), .C(n3979), .Y(n8111) );
  NAND2X1 U7635 ( .A(ram[3674]), .B(n12806), .Y(n3979) );
  OAI21X1 U7636 ( .A(n12713), .B(n12806), .C(n3980), .Y(n8112) );
  NAND2X1 U7637 ( .A(ram[3675]), .B(n12806), .Y(n3980) );
  OAI21X1 U7638 ( .A(n12707), .B(n12806), .C(n3981), .Y(n8113) );
  NAND2X1 U7639 ( .A(ram[3676]), .B(n12806), .Y(n3981) );
  OAI21X1 U7640 ( .A(n12701), .B(n12806), .C(n3982), .Y(n8114) );
  NAND2X1 U7641 ( .A(ram[3677]), .B(n12806), .Y(n3982) );
  OAI21X1 U7642 ( .A(n12695), .B(n12806), .C(n3983), .Y(n8115) );
  NAND2X1 U7643 ( .A(ram[3678]), .B(n12806), .Y(n3983) );
  OAI21X1 U7644 ( .A(n12689), .B(n12806), .C(n3984), .Y(n8116) );
  NAND2X1 U7645 ( .A(ram[3679]), .B(n12806), .Y(n3984) );
  OAI21X1 U7647 ( .A(n12779), .B(n12805), .C(n3986), .Y(n8117) );
  NAND2X1 U7648 ( .A(ram[3680]), .B(n12805), .Y(n3986) );
  OAI21X1 U7649 ( .A(n12773), .B(n12805), .C(n3987), .Y(n8118) );
  NAND2X1 U7650 ( .A(ram[3681]), .B(n12805), .Y(n3987) );
  OAI21X1 U7651 ( .A(n12767), .B(n12805), .C(n3988), .Y(n8119) );
  NAND2X1 U7652 ( .A(ram[3682]), .B(n12805), .Y(n3988) );
  OAI21X1 U7653 ( .A(n12761), .B(n12805), .C(n3989), .Y(n8120) );
  NAND2X1 U7654 ( .A(ram[3683]), .B(n12805), .Y(n3989) );
  OAI21X1 U7655 ( .A(n12755), .B(n12805), .C(n3990), .Y(n8121) );
  NAND2X1 U7656 ( .A(ram[3684]), .B(n12805), .Y(n3990) );
  OAI21X1 U7657 ( .A(n12749), .B(n12805), .C(n3991), .Y(n8122) );
  NAND2X1 U7658 ( .A(ram[3685]), .B(n12805), .Y(n3991) );
  OAI21X1 U7659 ( .A(n12743), .B(n12805), .C(n3992), .Y(n8123) );
  NAND2X1 U7660 ( .A(ram[3686]), .B(n12805), .Y(n3992) );
  OAI21X1 U7661 ( .A(n12737), .B(n12805), .C(n3993), .Y(n8124) );
  NAND2X1 U7662 ( .A(ram[3687]), .B(n12805), .Y(n3993) );
  OAI21X1 U7663 ( .A(n12731), .B(n12805), .C(n3994), .Y(n8125) );
  NAND2X1 U7664 ( .A(ram[3688]), .B(n12805), .Y(n3994) );
  OAI21X1 U7665 ( .A(n12725), .B(n12805), .C(n3995), .Y(n8126) );
  NAND2X1 U7666 ( .A(ram[3689]), .B(n12805), .Y(n3995) );
  OAI21X1 U7667 ( .A(n12719), .B(n12805), .C(n3996), .Y(n8127) );
  NAND2X1 U7668 ( .A(ram[3690]), .B(n12805), .Y(n3996) );
  OAI21X1 U7669 ( .A(n12713), .B(n12805), .C(n3997), .Y(n8128) );
  NAND2X1 U7670 ( .A(ram[3691]), .B(n12805), .Y(n3997) );
  OAI21X1 U7671 ( .A(n12707), .B(n12805), .C(n3998), .Y(n8129) );
  NAND2X1 U7672 ( .A(ram[3692]), .B(n12805), .Y(n3998) );
  OAI21X1 U7673 ( .A(n12701), .B(n12805), .C(n3999), .Y(n8130) );
  NAND2X1 U7674 ( .A(ram[3693]), .B(n12805), .Y(n3999) );
  OAI21X1 U7675 ( .A(n12695), .B(n12805), .C(n4000), .Y(n8131) );
  NAND2X1 U7676 ( .A(ram[3694]), .B(n12805), .Y(n4000) );
  OAI21X1 U7677 ( .A(n12689), .B(n12805), .C(n4001), .Y(n8132) );
  NAND2X1 U7678 ( .A(ram[3695]), .B(n12805), .Y(n4001) );
  OAI21X1 U7680 ( .A(n12779), .B(n12804), .C(n4003), .Y(n8133) );
  NAND2X1 U7681 ( .A(ram[3696]), .B(n12804), .Y(n4003) );
  OAI21X1 U7682 ( .A(n12773), .B(n12804), .C(n4004), .Y(n8134) );
  NAND2X1 U7683 ( .A(ram[3697]), .B(n12804), .Y(n4004) );
  OAI21X1 U7684 ( .A(n12767), .B(n12804), .C(n4005), .Y(n8135) );
  NAND2X1 U7685 ( .A(ram[3698]), .B(n12804), .Y(n4005) );
  OAI21X1 U7686 ( .A(n12761), .B(n12804), .C(n4006), .Y(n8136) );
  NAND2X1 U7687 ( .A(ram[3699]), .B(n12804), .Y(n4006) );
  OAI21X1 U7688 ( .A(n12755), .B(n12804), .C(n4007), .Y(n8137) );
  NAND2X1 U7689 ( .A(ram[3700]), .B(n12804), .Y(n4007) );
  OAI21X1 U7690 ( .A(n12749), .B(n12804), .C(n4008), .Y(n8138) );
  NAND2X1 U7691 ( .A(ram[3701]), .B(n12804), .Y(n4008) );
  OAI21X1 U7692 ( .A(n12743), .B(n12804), .C(n4009), .Y(n8139) );
  NAND2X1 U7693 ( .A(ram[3702]), .B(n12804), .Y(n4009) );
  OAI21X1 U7694 ( .A(n12737), .B(n12804), .C(n4010), .Y(n8140) );
  NAND2X1 U7695 ( .A(ram[3703]), .B(n12804), .Y(n4010) );
  OAI21X1 U7696 ( .A(n12731), .B(n12804), .C(n4011), .Y(n8141) );
  NAND2X1 U7697 ( .A(ram[3704]), .B(n12804), .Y(n4011) );
  OAI21X1 U7698 ( .A(n12725), .B(n12804), .C(n4012), .Y(n8142) );
  NAND2X1 U7699 ( .A(ram[3705]), .B(n12804), .Y(n4012) );
  OAI21X1 U7700 ( .A(n12719), .B(n12804), .C(n4013), .Y(n8143) );
  NAND2X1 U7701 ( .A(ram[3706]), .B(n12804), .Y(n4013) );
  OAI21X1 U7702 ( .A(n12713), .B(n12804), .C(n4014), .Y(n8144) );
  NAND2X1 U7703 ( .A(ram[3707]), .B(n12804), .Y(n4014) );
  OAI21X1 U7704 ( .A(n12707), .B(n12804), .C(n4015), .Y(n8145) );
  NAND2X1 U7705 ( .A(ram[3708]), .B(n12804), .Y(n4015) );
  OAI21X1 U7706 ( .A(n12701), .B(n12804), .C(n4016), .Y(n8146) );
  NAND2X1 U7707 ( .A(ram[3709]), .B(n12804), .Y(n4016) );
  OAI21X1 U7708 ( .A(n12695), .B(n12804), .C(n4017), .Y(n8147) );
  NAND2X1 U7709 ( .A(ram[3710]), .B(n12804), .Y(n4017) );
  OAI21X1 U7710 ( .A(n12689), .B(n12804), .C(n4018), .Y(n8148) );
  NAND2X1 U7711 ( .A(ram[3711]), .B(n12804), .Y(n4018) );
  OAI21X1 U7713 ( .A(n12779), .B(n12803), .C(n4020), .Y(n8149) );
  NAND2X1 U7714 ( .A(ram[3712]), .B(n12803), .Y(n4020) );
  OAI21X1 U7715 ( .A(n12773), .B(n12803), .C(n4021), .Y(n8150) );
  NAND2X1 U7716 ( .A(ram[3713]), .B(n12803), .Y(n4021) );
  OAI21X1 U7717 ( .A(n12767), .B(n12803), .C(n4022), .Y(n8151) );
  NAND2X1 U7718 ( .A(ram[3714]), .B(n12803), .Y(n4022) );
  OAI21X1 U7719 ( .A(n12761), .B(n12803), .C(n4023), .Y(n8152) );
  NAND2X1 U7720 ( .A(ram[3715]), .B(n12803), .Y(n4023) );
  OAI21X1 U7721 ( .A(n12755), .B(n12803), .C(n4024), .Y(n8153) );
  NAND2X1 U7722 ( .A(ram[3716]), .B(n12803), .Y(n4024) );
  OAI21X1 U7723 ( .A(n12749), .B(n12803), .C(n4025), .Y(n8154) );
  NAND2X1 U7724 ( .A(ram[3717]), .B(n12803), .Y(n4025) );
  OAI21X1 U7725 ( .A(n12743), .B(n12803), .C(n4026), .Y(n8155) );
  NAND2X1 U7726 ( .A(ram[3718]), .B(n12803), .Y(n4026) );
  OAI21X1 U7727 ( .A(n12737), .B(n12803), .C(n4027), .Y(n8156) );
  NAND2X1 U7728 ( .A(ram[3719]), .B(n12803), .Y(n4027) );
  OAI21X1 U7729 ( .A(n12731), .B(n12803), .C(n4028), .Y(n8157) );
  NAND2X1 U7730 ( .A(ram[3720]), .B(n12803), .Y(n4028) );
  OAI21X1 U7731 ( .A(n12725), .B(n12803), .C(n4029), .Y(n8158) );
  NAND2X1 U7732 ( .A(ram[3721]), .B(n12803), .Y(n4029) );
  OAI21X1 U7733 ( .A(n12719), .B(n12803), .C(n4030), .Y(n8159) );
  NAND2X1 U7734 ( .A(ram[3722]), .B(n12803), .Y(n4030) );
  OAI21X1 U7735 ( .A(n12713), .B(n12803), .C(n4031), .Y(n8160) );
  NAND2X1 U7736 ( .A(ram[3723]), .B(n12803), .Y(n4031) );
  OAI21X1 U7737 ( .A(n12707), .B(n12803), .C(n4032), .Y(n8161) );
  NAND2X1 U7738 ( .A(ram[3724]), .B(n12803), .Y(n4032) );
  OAI21X1 U7739 ( .A(n12701), .B(n12803), .C(n4033), .Y(n8162) );
  NAND2X1 U7740 ( .A(ram[3725]), .B(n12803), .Y(n4033) );
  OAI21X1 U7741 ( .A(n12695), .B(n12803), .C(n4034), .Y(n8163) );
  NAND2X1 U7742 ( .A(ram[3726]), .B(n12803), .Y(n4034) );
  OAI21X1 U7743 ( .A(n12689), .B(n12803), .C(n4035), .Y(n8164) );
  NAND2X1 U7744 ( .A(ram[3727]), .B(n12803), .Y(n4035) );
  OAI21X1 U7746 ( .A(n12779), .B(n12802), .C(n4037), .Y(n8165) );
  NAND2X1 U7747 ( .A(ram[3728]), .B(n12802), .Y(n4037) );
  OAI21X1 U7748 ( .A(n12773), .B(n12802), .C(n4038), .Y(n8166) );
  NAND2X1 U7749 ( .A(ram[3729]), .B(n12802), .Y(n4038) );
  OAI21X1 U7750 ( .A(n12767), .B(n12802), .C(n4039), .Y(n8167) );
  NAND2X1 U7751 ( .A(ram[3730]), .B(n12802), .Y(n4039) );
  OAI21X1 U7752 ( .A(n12761), .B(n12802), .C(n4040), .Y(n8168) );
  NAND2X1 U7753 ( .A(ram[3731]), .B(n12802), .Y(n4040) );
  OAI21X1 U7754 ( .A(n12755), .B(n12802), .C(n4041), .Y(n8169) );
  NAND2X1 U7755 ( .A(ram[3732]), .B(n12802), .Y(n4041) );
  OAI21X1 U7756 ( .A(n12749), .B(n12802), .C(n4042), .Y(n8170) );
  NAND2X1 U7757 ( .A(ram[3733]), .B(n12802), .Y(n4042) );
  OAI21X1 U7758 ( .A(n12743), .B(n12802), .C(n4043), .Y(n8171) );
  NAND2X1 U7759 ( .A(ram[3734]), .B(n12802), .Y(n4043) );
  OAI21X1 U7760 ( .A(n12737), .B(n12802), .C(n4044), .Y(n8172) );
  NAND2X1 U7761 ( .A(ram[3735]), .B(n12802), .Y(n4044) );
  OAI21X1 U7762 ( .A(n12731), .B(n12802), .C(n4045), .Y(n8173) );
  NAND2X1 U7763 ( .A(ram[3736]), .B(n12802), .Y(n4045) );
  OAI21X1 U7764 ( .A(n12725), .B(n12802), .C(n4046), .Y(n8174) );
  NAND2X1 U7765 ( .A(ram[3737]), .B(n12802), .Y(n4046) );
  OAI21X1 U7766 ( .A(n12719), .B(n12802), .C(n4047), .Y(n8175) );
  NAND2X1 U7767 ( .A(ram[3738]), .B(n12802), .Y(n4047) );
  OAI21X1 U7768 ( .A(n12713), .B(n12802), .C(n4048), .Y(n8176) );
  NAND2X1 U7769 ( .A(ram[3739]), .B(n12802), .Y(n4048) );
  OAI21X1 U7770 ( .A(n12707), .B(n12802), .C(n4049), .Y(n8177) );
  NAND2X1 U7771 ( .A(ram[3740]), .B(n12802), .Y(n4049) );
  OAI21X1 U7772 ( .A(n12701), .B(n12802), .C(n4050), .Y(n8178) );
  NAND2X1 U7773 ( .A(ram[3741]), .B(n12802), .Y(n4050) );
  OAI21X1 U7774 ( .A(n12695), .B(n12802), .C(n4051), .Y(n8179) );
  NAND2X1 U7775 ( .A(ram[3742]), .B(n12802), .Y(n4051) );
  OAI21X1 U7776 ( .A(n12689), .B(n12802), .C(n4052), .Y(n8180) );
  NAND2X1 U7777 ( .A(ram[3743]), .B(n12802), .Y(n4052) );
  OAI21X1 U7779 ( .A(n12779), .B(n12801), .C(n4054), .Y(n8181) );
  NAND2X1 U7780 ( .A(ram[3744]), .B(n12801), .Y(n4054) );
  OAI21X1 U7781 ( .A(n12773), .B(n12801), .C(n4055), .Y(n8182) );
  NAND2X1 U7782 ( .A(ram[3745]), .B(n12801), .Y(n4055) );
  OAI21X1 U7783 ( .A(n12767), .B(n12801), .C(n4056), .Y(n8183) );
  NAND2X1 U7784 ( .A(ram[3746]), .B(n12801), .Y(n4056) );
  OAI21X1 U7785 ( .A(n12761), .B(n12801), .C(n4057), .Y(n8184) );
  NAND2X1 U7786 ( .A(ram[3747]), .B(n12801), .Y(n4057) );
  OAI21X1 U7787 ( .A(n12755), .B(n12801), .C(n4058), .Y(n8185) );
  NAND2X1 U7788 ( .A(ram[3748]), .B(n12801), .Y(n4058) );
  OAI21X1 U7789 ( .A(n12749), .B(n12801), .C(n4059), .Y(n8186) );
  NAND2X1 U7790 ( .A(ram[3749]), .B(n12801), .Y(n4059) );
  OAI21X1 U7791 ( .A(n12743), .B(n12801), .C(n4060), .Y(n8187) );
  NAND2X1 U7792 ( .A(ram[3750]), .B(n12801), .Y(n4060) );
  OAI21X1 U7793 ( .A(n12737), .B(n12801), .C(n4061), .Y(n8188) );
  NAND2X1 U7794 ( .A(ram[3751]), .B(n12801), .Y(n4061) );
  OAI21X1 U7795 ( .A(n12731), .B(n12801), .C(n4062), .Y(n8189) );
  NAND2X1 U7796 ( .A(ram[3752]), .B(n12801), .Y(n4062) );
  OAI21X1 U7797 ( .A(n12725), .B(n12801), .C(n4063), .Y(n8190) );
  NAND2X1 U7798 ( .A(ram[3753]), .B(n12801), .Y(n4063) );
  OAI21X1 U7799 ( .A(n12719), .B(n12801), .C(n4064), .Y(n8191) );
  NAND2X1 U7800 ( .A(ram[3754]), .B(n12801), .Y(n4064) );
  OAI21X1 U7801 ( .A(n12713), .B(n12801), .C(n4065), .Y(n8192) );
  NAND2X1 U7802 ( .A(ram[3755]), .B(n12801), .Y(n4065) );
  OAI21X1 U7803 ( .A(n12707), .B(n12801), .C(n4066), .Y(n8193) );
  NAND2X1 U7804 ( .A(ram[3756]), .B(n12801), .Y(n4066) );
  OAI21X1 U7805 ( .A(n12701), .B(n12801), .C(n4067), .Y(n8194) );
  NAND2X1 U7806 ( .A(ram[3757]), .B(n12801), .Y(n4067) );
  OAI21X1 U7807 ( .A(n12695), .B(n12801), .C(n4068), .Y(n8195) );
  NAND2X1 U7808 ( .A(ram[3758]), .B(n12801), .Y(n4068) );
  OAI21X1 U7809 ( .A(n12689), .B(n12801), .C(n4069), .Y(n8196) );
  NAND2X1 U7810 ( .A(ram[3759]), .B(n12801), .Y(n4069) );
  OAI21X1 U7812 ( .A(n12778), .B(n12800), .C(n4071), .Y(n8197) );
  NAND2X1 U7813 ( .A(ram[3760]), .B(n12800), .Y(n4071) );
  OAI21X1 U7814 ( .A(n12772), .B(n12800), .C(n4072), .Y(n8198) );
  NAND2X1 U7815 ( .A(ram[3761]), .B(n12800), .Y(n4072) );
  OAI21X1 U7816 ( .A(n12766), .B(n12800), .C(n4073), .Y(n8199) );
  NAND2X1 U7817 ( .A(ram[3762]), .B(n12800), .Y(n4073) );
  OAI21X1 U7818 ( .A(n12760), .B(n12800), .C(n4074), .Y(n8200) );
  NAND2X1 U7819 ( .A(ram[3763]), .B(n12800), .Y(n4074) );
  OAI21X1 U7820 ( .A(n12754), .B(n12800), .C(n4075), .Y(n8201) );
  NAND2X1 U7821 ( .A(ram[3764]), .B(n12800), .Y(n4075) );
  OAI21X1 U7822 ( .A(n12748), .B(n12800), .C(n4076), .Y(n8202) );
  NAND2X1 U7823 ( .A(ram[3765]), .B(n12800), .Y(n4076) );
  OAI21X1 U7824 ( .A(n12742), .B(n12800), .C(n4077), .Y(n8203) );
  NAND2X1 U7825 ( .A(ram[3766]), .B(n12800), .Y(n4077) );
  OAI21X1 U7826 ( .A(n12736), .B(n12800), .C(n4078), .Y(n8204) );
  NAND2X1 U7827 ( .A(ram[3767]), .B(n12800), .Y(n4078) );
  OAI21X1 U7828 ( .A(n12730), .B(n12800), .C(n4079), .Y(n8205) );
  NAND2X1 U7829 ( .A(ram[3768]), .B(n12800), .Y(n4079) );
  OAI21X1 U7830 ( .A(n12724), .B(n12800), .C(n4080), .Y(n8206) );
  NAND2X1 U7831 ( .A(ram[3769]), .B(n12800), .Y(n4080) );
  OAI21X1 U7832 ( .A(n12718), .B(n12800), .C(n4081), .Y(n8207) );
  NAND2X1 U7833 ( .A(ram[3770]), .B(n12800), .Y(n4081) );
  OAI21X1 U7834 ( .A(n12712), .B(n12800), .C(n4082), .Y(n8208) );
  NAND2X1 U7835 ( .A(ram[3771]), .B(n12800), .Y(n4082) );
  OAI21X1 U7836 ( .A(n12706), .B(n12800), .C(n4083), .Y(n8209) );
  NAND2X1 U7837 ( .A(ram[3772]), .B(n12800), .Y(n4083) );
  OAI21X1 U7838 ( .A(n12700), .B(n12800), .C(n4084), .Y(n8210) );
  NAND2X1 U7839 ( .A(ram[3773]), .B(n12800), .Y(n4084) );
  OAI21X1 U7840 ( .A(n12694), .B(n12800), .C(n4085), .Y(n8211) );
  NAND2X1 U7841 ( .A(ram[3774]), .B(n12800), .Y(n4085) );
  OAI21X1 U7842 ( .A(n12688), .B(n12800), .C(n4086), .Y(n8212) );
  NAND2X1 U7843 ( .A(ram[3775]), .B(n12800), .Y(n4086) );
  OAI21X1 U7845 ( .A(n12777), .B(n12799), .C(n4088), .Y(n8213) );
  NAND2X1 U7846 ( .A(ram[3776]), .B(n12799), .Y(n4088) );
  OAI21X1 U7847 ( .A(n12771), .B(n12799), .C(n4089), .Y(n8214) );
  NAND2X1 U7848 ( .A(ram[3777]), .B(n12799), .Y(n4089) );
  OAI21X1 U7849 ( .A(n12765), .B(n12799), .C(n4090), .Y(n8215) );
  NAND2X1 U7850 ( .A(ram[3778]), .B(n12799), .Y(n4090) );
  OAI21X1 U7851 ( .A(n12759), .B(n12799), .C(n4091), .Y(n8216) );
  NAND2X1 U7852 ( .A(ram[3779]), .B(n12799), .Y(n4091) );
  OAI21X1 U7853 ( .A(n12753), .B(n12799), .C(n4092), .Y(n8217) );
  NAND2X1 U7854 ( .A(ram[3780]), .B(n12799), .Y(n4092) );
  OAI21X1 U7855 ( .A(n12747), .B(n12799), .C(n4093), .Y(n8218) );
  NAND2X1 U7856 ( .A(ram[3781]), .B(n12799), .Y(n4093) );
  OAI21X1 U7857 ( .A(n12741), .B(n12799), .C(n4094), .Y(n8219) );
  NAND2X1 U7858 ( .A(ram[3782]), .B(n12799), .Y(n4094) );
  OAI21X1 U7859 ( .A(n12735), .B(n12799), .C(n4095), .Y(n8220) );
  NAND2X1 U7860 ( .A(ram[3783]), .B(n12799), .Y(n4095) );
  OAI21X1 U7861 ( .A(n12729), .B(n12799), .C(n4096), .Y(n8221) );
  NAND2X1 U7862 ( .A(ram[3784]), .B(n12799), .Y(n4096) );
  OAI21X1 U7863 ( .A(n12723), .B(n12799), .C(n4097), .Y(n8222) );
  NAND2X1 U7864 ( .A(ram[3785]), .B(n12799), .Y(n4097) );
  OAI21X1 U7865 ( .A(n12717), .B(n12799), .C(n4098), .Y(n8223) );
  NAND2X1 U7866 ( .A(ram[3786]), .B(n12799), .Y(n4098) );
  OAI21X1 U7867 ( .A(n12711), .B(n12799), .C(n4099), .Y(n8224) );
  NAND2X1 U7868 ( .A(ram[3787]), .B(n12799), .Y(n4099) );
  OAI21X1 U7869 ( .A(n12705), .B(n12799), .C(n4100), .Y(n8225) );
  NAND2X1 U7870 ( .A(ram[3788]), .B(n12799), .Y(n4100) );
  OAI21X1 U7871 ( .A(n12699), .B(n12799), .C(n4101), .Y(n8226) );
  NAND2X1 U7872 ( .A(ram[3789]), .B(n12799), .Y(n4101) );
  OAI21X1 U7873 ( .A(n12693), .B(n12799), .C(n4102), .Y(n8227) );
  NAND2X1 U7874 ( .A(ram[3790]), .B(n12799), .Y(n4102) );
  OAI21X1 U7875 ( .A(n12687), .B(n12799), .C(n4103), .Y(n8228) );
  NAND2X1 U7876 ( .A(ram[3791]), .B(n12799), .Y(n4103) );
  OAI21X1 U7878 ( .A(n12776), .B(n12798), .C(n4105), .Y(n8229) );
  NAND2X1 U7879 ( .A(ram[3792]), .B(n12798), .Y(n4105) );
  OAI21X1 U7880 ( .A(n12770), .B(n12798), .C(n4106), .Y(n8230) );
  NAND2X1 U7881 ( .A(ram[3793]), .B(n12798), .Y(n4106) );
  OAI21X1 U7882 ( .A(n12764), .B(n12798), .C(n4107), .Y(n8231) );
  NAND2X1 U7883 ( .A(ram[3794]), .B(n12798), .Y(n4107) );
  OAI21X1 U7884 ( .A(n12758), .B(n12798), .C(n4108), .Y(n8232) );
  NAND2X1 U7885 ( .A(ram[3795]), .B(n12798), .Y(n4108) );
  OAI21X1 U7886 ( .A(n12752), .B(n12798), .C(n4109), .Y(n8233) );
  NAND2X1 U7887 ( .A(ram[3796]), .B(n12798), .Y(n4109) );
  OAI21X1 U7888 ( .A(n12746), .B(n12798), .C(n4110), .Y(n8234) );
  NAND2X1 U7889 ( .A(ram[3797]), .B(n12798), .Y(n4110) );
  OAI21X1 U7890 ( .A(n12740), .B(n12798), .C(n4111), .Y(n8235) );
  NAND2X1 U7891 ( .A(ram[3798]), .B(n12798), .Y(n4111) );
  OAI21X1 U7892 ( .A(n12734), .B(n12798), .C(n4112), .Y(n8236) );
  NAND2X1 U7893 ( .A(ram[3799]), .B(n12798), .Y(n4112) );
  OAI21X1 U7894 ( .A(n12728), .B(n12798), .C(n4113), .Y(n8237) );
  NAND2X1 U7895 ( .A(ram[3800]), .B(n12798), .Y(n4113) );
  OAI21X1 U7896 ( .A(n12722), .B(n12798), .C(n4114), .Y(n8238) );
  NAND2X1 U7897 ( .A(ram[3801]), .B(n12798), .Y(n4114) );
  OAI21X1 U7898 ( .A(n12716), .B(n12798), .C(n4115), .Y(n8239) );
  NAND2X1 U7899 ( .A(ram[3802]), .B(n12798), .Y(n4115) );
  OAI21X1 U7900 ( .A(n12710), .B(n12798), .C(n4116), .Y(n8240) );
  NAND2X1 U7901 ( .A(ram[3803]), .B(n12798), .Y(n4116) );
  OAI21X1 U7902 ( .A(n12704), .B(n12798), .C(n4117), .Y(n8241) );
  NAND2X1 U7903 ( .A(ram[3804]), .B(n12798), .Y(n4117) );
  OAI21X1 U7904 ( .A(n12698), .B(n12798), .C(n4118), .Y(n8242) );
  NAND2X1 U7905 ( .A(ram[3805]), .B(n12798), .Y(n4118) );
  OAI21X1 U7906 ( .A(n12692), .B(n12798), .C(n4119), .Y(n8243) );
  NAND2X1 U7907 ( .A(ram[3806]), .B(n12798), .Y(n4119) );
  OAI21X1 U7908 ( .A(n12686), .B(n12798), .C(n4120), .Y(n8244) );
  NAND2X1 U7909 ( .A(ram[3807]), .B(n12798), .Y(n4120) );
  OAI21X1 U7911 ( .A(n12779), .B(n12797), .C(n4122), .Y(n8245) );
  NAND2X1 U7912 ( .A(ram[3808]), .B(n12797), .Y(n4122) );
  OAI21X1 U7913 ( .A(n12773), .B(n12797), .C(n4123), .Y(n8246) );
  NAND2X1 U7914 ( .A(ram[3809]), .B(n12797), .Y(n4123) );
  OAI21X1 U7915 ( .A(n12767), .B(n12797), .C(n4124), .Y(n8247) );
  NAND2X1 U7916 ( .A(ram[3810]), .B(n12797), .Y(n4124) );
  OAI21X1 U7917 ( .A(n12761), .B(n12797), .C(n4125), .Y(n8248) );
  NAND2X1 U7918 ( .A(ram[3811]), .B(n12797), .Y(n4125) );
  OAI21X1 U7919 ( .A(n12755), .B(n12797), .C(n4126), .Y(n8249) );
  NAND2X1 U7920 ( .A(ram[3812]), .B(n12797), .Y(n4126) );
  OAI21X1 U7921 ( .A(n12749), .B(n12797), .C(n4127), .Y(n8250) );
  NAND2X1 U7922 ( .A(ram[3813]), .B(n12797), .Y(n4127) );
  OAI21X1 U7923 ( .A(n12743), .B(n12797), .C(n4128), .Y(n8251) );
  NAND2X1 U7924 ( .A(ram[3814]), .B(n12797), .Y(n4128) );
  OAI21X1 U7925 ( .A(n12737), .B(n12797), .C(n4129), .Y(n8252) );
  NAND2X1 U7926 ( .A(ram[3815]), .B(n12797), .Y(n4129) );
  OAI21X1 U7927 ( .A(n12731), .B(n12797), .C(n4130), .Y(n8253) );
  NAND2X1 U7928 ( .A(ram[3816]), .B(n12797), .Y(n4130) );
  OAI21X1 U7929 ( .A(n12725), .B(n12797), .C(n4131), .Y(n8254) );
  NAND2X1 U7930 ( .A(ram[3817]), .B(n12797), .Y(n4131) );
  OAI21X1 U7931 ( .A(n12719), .B(n12797), .C(n4132), .Y(n8255) );
  NAND2X1 U7932 ( .A(ram[3818]), .B(n12797), .Y(n4132) );
  OAI21X1 U7933 ( .A(n12713), .B(n12797), .C(n4133), .Y(n8256) );
  NAND2X1 U7934 ( .A(ram[3819]), .B(n12797), .Y(n4133) );
  OAI21X1 U7935 ( .A(n12707), .B(n12797), .C(n4134), .Y(n8257) );
  NAND2X1 U7936 ( .A(ram[3820]), .B(n12797), .Y(n4134) );
  OAI21X1 U7937 ( .A(n12701), .B(n12797), .C(n4135), .Y(n8258) );
  NAND2X1 U7938 ( .A(ram[3821]), .B(n12797), .Y(n4135) );
  OAI21X1 U7939 ( .A(n12695), .B(n12797), .C(n4136), .Y(n8259) );
  NAND2X1 U7940 ( .A(ram[3822]), .B(n12797), .Y(n4136) );
  OAI21X1 U7941 ( .A(n12689), .B(n12797), .C(n4137), .Y(n8260) );
  NAND2X1 U7942 ( .A(ram[3823]), .B(n12797), .Y(n4137) );
  OAI21X1 U7944 ( .A(n12778), .B(n12796), .C(n4139), .Y(n8261) );
  NAND2X1 U7945 ( .A(ram[3824]), .B(n12796), .Y(n4139) );
  OAI21X1 U7946 ( .A(n12772), .B(n12796), .C(n4140), .Y(n8262) );
  NAND2X1 U7947 ( .A(ram[3825]), .B(n12796), .Y(n4140) );
  OAI21X1 U7948 ( .A(n12766), .B(n12796), .C(n4141), .Y(n8263) );
  NAND2X1 U7949 ( .A(ram[3826]), .B(n12796), .Y(n4141) );
  OAI21X1 U7950 ( .A(n12760), .B(n12796), .C(n4142), .Y(n8264) );
  NAND2X1 U7951 ( .A(ram[3827]), .B(n12796), .Y(n4142) );
  OAI21X1 U7952 ( .A(n12754), .B(n12796), .C(n4143), .Y(n8265) );
  NAND2X1 U7953 ( .A(ram[3828]), .B(n12796), .Y(n4143) );
  OAI21X1 U7954 ( .A(n12748), .B(n12796), .C(n4144), .Y(n8266) );
  NAND2X1 U7955 ( .A(ram[3829]), .B(n12796), .Y(n4144) );
  OAI21X1 U7956 ( .A(n12742), .B(n12796), .C(n4145), .Y(n8267) );
  NAND2X1 U7957 ( .A(ram[3830]), .B(n12796), .Y(n4145) );
  OAI21X1 U7958 ( .A(n12736), .B(n12796), .C(n4146), .Y(n8268) );
  NAND2X1 U7959 ( .A(ram[3831]), .B(n12796), .Y(n4146) );
  OAI21X1 U7960 ( .A(n12730), .B(n12796), .C(n4147), .Y(n8269) );
  NAND2X1 U7961 ( .A(ram[3832]), .B(n12796), .Y(n4147) );
  OAI21X1 U7962 ( .A(n12724), .B(n12796), .C(n4148), .Y(n8270) );
  NAND2X1 U7963 ( .A(ram[3833]), .B(n12796), .Y(n4148) );
  OAI21X1 U7964 ( .A(n12718), .B(n12796), .C(n4149), .Y(n8271) );
  NAND2X1 U7965 ( .A(ram[3834]), .B(n12796), .Y(n4149) );
  OAI21X1 U7966 ( .A(n12712), .B(n12796), .C(n4150), .Y(n8272) );
  NAND2X1 U7967 ( .A(ram[3835]), .B(n12796), .Y(n4150) );
  OAI21X1 U7968 ( .A(n12706), .B(n12796), .C(n4151), .Y(n8273) );
  NAND2X1 U7969 ( .A(ram[3836]), .B(n12796), .Y(n4151) );
  OAI21X1 U7970 ( .A(n12700), .B(n12796), .C(n4152), .Y(n8274) );
  NAND2X1 U7971 ( .A(ram[3837]), .B(n12796), .Y(n4152) );
  OAI21X1 U7972 ( .A(n12694), .B(n12796), .C(n4153), .Y(n8275) );
  NAND2X1 U7973 ( .A(ram[3838]), .B(n12796), .Y(n4153) );
  OAI21X1 U7974 ( .A(n12688), .B(n12796), .C(n4154), .Y(n8276) );
  NAND2X1 U7975 ( .A(ram[3839]), .B(n12796), .Y(n4154) );
  NAND3X1 U7977 ( .A(n875), .B(mem_write_en), .C(n3609), .Y(n4155) );
  AND2X1 U7978 ( .A(mem_access_addr[5]), .B(n13038), .Y(n875) );
  OAI21X1 U7979 ( .A(n12777), .B(n12795), .C(n4157), .Y(n8277) );
  NAND2X1 U7980 ( .A(ram[3840]), .B(n12795), .Y(n4157) );
  OAI21X1 U7981 ( .A(n12771), .B(n12795), .C(n4158), .Y(n8278) );
  NAND2X1 U7982 ( .A(ram[3841]), .B(n12795), .Y(n4158) );
  OAI21X1 U7983 ( .A(n12765), .B(n12795), .C(n4159), .Y(n8279) );
  NAND2X1 U7984 ( .A(ram[3842]), .B(n12795), .Y(n4159) );
  OAI21X1 U7985 ( .A(n12759), .B(n12795), .C(n4160), .Y(n8280) );
  NAND2X1 U7986 ( .A(ram[3843]), .B(n12795), .Y(n4160) );
  OAI21X1 U7987 ( .A(n12753), .B(n12795), .C(n4161), .Y(n8281) );
  NAND2X1 U7988 ( .A(ram[3844]), .B(n12795), .Y(n4161) );
  OAI21X1 U7989 ( .A(n12747), .B(n12795), .C(n4162), .Y(n8282) );
  NAND2X1 U7990 ( .A(ram[3845]), .B(n12795), .Y(n4162) );
  OAI21X1 U7991 ( .A(n12741), .B(n12795), .C(n4163), .Y(n8283) );
  NAND2X1 U7992 ( .A(ram[3846]), .B(n12795), .Y(n4163) );
  OAI21X1 U7993 ( .A(n12735), .B(n12795), .C(n4164), .Y(n8284) );
  NAND2X1 U7994 ( .A(ram[3847]), .B(n12795), .Y(n4164) );
  OAI21X1 U7995 ( .A(n12729), .B(n12795), .C(n4165), .Y(n8285) );
  NAND2X1 U7996 ( .A(ram[3848]), .B(n12795), .Y(n4165) );
  OAI21X1 U7997 ( .A(n12723), .B(n12795), .C(n4166), .Y(n8286) );
  NAND2X1 U7998 ( .A(ram[3849]), .B(n12795), .Y(n4166) );
  OAI21X1 U7999 ( .A(n12717), .B(n12795), .C(n4167), .Y(n8287) );
  NAND2X1 U8000 ( .A(ram[3850]), .B(n12795), .Y(n4167) );
  OAI21X1 U8001 ( .A(n12711), .B(n12795), .C(n4168), .Y(n8288) );
  NAND2X1 U8002 ( .A(ram[3851]), .B(n12795), .Y(n4168) );
  OAI21X1 U8003 ( .A(n12705), .B(n12795), .C(n4169), .Y(n8289) );
  NAND2X1 U8004 ( .A(ram[3852]), .B(n12795), .Y(n4169) );
  OAI21X1 U8005 ( .A(n12699), .B(n12795), .C(n4170), .Y(n8290) );
  NAND2X1 U8006 ( .A(ram[3853]), .B(n12795), .Y(n4170) );
  OAI21X1 U8007 ( .A(n12693), .B(n12795), .C(n4171), .Y(n8291) );
  NAND2X1 U8008 ( .A(ram[3854]), .B(n12795), .Y(n4171) );
  OAI21X1 U8009 ( .A(n12687), .B(n12795), .C(n4172), .Y(n8292) );
  NAND2X1 U8010 ( .A(ram[3855]), .B(n12795), .Y(n4172) );
  OAI21X1 U8013 ( .A(n12776), .B(n12794), .C(n4176), .Y(n8293) );
  NAND2X1 U8014 ( .A(ram[3856]), .B(n12794), .Y(n4176) );
  OAI21X1 U8015 ( .A(n12770), .B(n12794), .C(n4177), .Y(n8294) );
  NAND2X1 U8016 ( .A(ram[3857]), .B(n12794), .Y(n4177) );
  OAI21X1 U8017 ( .A(n12764), .B(n12794), .C(n4178), .Y(n8295) );
  NAND2X1 U8018 ( .A(ram[3858]), .B(n12794), .Y(n4178) );
  OAI21X1 U8019 ( .A(n12758), .B(n12794), .C(n4179), .Y(n8296) );
  NAND2X1 U8020 ( .A(ram[3859]), .B(n12794), .Y(n4179) );
  OAI21X1 U8021 ( .A(n12752), .B(n12794), .C(n4180), .Y(n8297) );
  NAND2X1 U8022 ( .A(ram[3860]), .B(n12794), .Y(n4180) );
  OAI21X1 U8023 ( .A(n12746), .B(n12794), .C(n4181), .Y(n8298) );
  NAND2X1 U8024 ( .A(ram[3861]), .B(n12794), .Y(n4181) );
  OAI21X1 U8025 ( .A(n12740), .B(n12794), .C(n4182), .Y(n8299) );
  NAND2X1 U8026 ( .A(ram[3862]), .B(n12794), .Y(n4182) );
  OAI21X1 U8027 ( .A(n12734), .B(n12794), .C(n4183), .Y(n8300) );
  NAND2X1 U8028 ( .A(ram[3863]), .B(n12794), .Y(n4183) );
  OAI21X1 U8029 ( .A(n12728), .B(n12794), .C(n4184), .Y(n8301) );
  NAND2X1 U8030 ( .A(ram[3864]), .B(n12794), .Y(n4184) );
  OAI21X1 U8031 ( .A(n12722), .B(n12794), .C(n4185), .Y(n8302) );
  NAND2X1 U8032 ( .A(ram[3865]), .B(n12794), .Y(n4185) );
  OAI21X1 U8033 ( .A(n12716), .B(n12794), .C(n4186), .Y(n8303) );
  NAND2X1 U8034 ( .A(ram[3866]), .B(n12794), .Y(n4186) );
  OAI21X1 U8035 ( .A(n12710), .B(n12794), .C(n4187), .Y(n8304) );
  NAND2X1 U8036 ( .A(ram[3867]), .B(n12794), .Y(n4187) );
  OAI21X1 U8037 ( .A(n12704), .B(n12794), .C(n4188), .Y(n8305) );
  NAND2X1 U8038 ( .A(ram[3868]), .B(n12794), .Y(n4188) );
  OAI21X1 U8039 ( .A(n12698), .B(n12794), .C(n4189), .Y(n8306) );
  NAND2X1 U8040 ( .A(ram[3869]), .B(n12794), .Y(n4189) );
  OAI21X1 U8041 ( .A(n12692), .B(n12794), .C(n4190), .Y(n8307) );
  NAND2X1 U8042 ( .A(ram[3870]), .B(n12794), .Y(n4190) );
  OAI21X1 U8043 ( .A(n12686), .B(n12794), .C(n4191), .Y(n8308) );
  NAND2X1 U8044 ( .A(ram[3871]), .B(n12794), .Y(n4191) );
  OAI21X1 U8047 ( .A(n12779), .B(n12793), .C(n4194), .Y(n8309) );
  NAND2X1 U8048 ( .A(ram[3872]), .B(n12793), .Y(n4194) );
  OAI21X1 U8049 ( .A(n12773), .B(n12793), .C(n4195), .Y(n8310) );
  NAND2X1 U8050 ( .A(ram[3873]), .B(n12793), .Y(n4195) );
  OAI21X1 U8051 ( .A(n12767), .B(n12793), .C(n4196), .Y(n8311) );
  NAND2X1 U8052 ( .A(ram[3874]), .B(n12793), .Y(n4196) );
  OAI21X1 U8053 ( .A(n12761), .B(n12793), .C(n4197), .Y(n8312) );
  NAND2X1 U8054 ( .A(ram[3875]), .B(n12793), .Y(n4197) );
  OAI21X1 U8055 ( .A(n12755), .B(n12793), .C(n4198), .Y(n8313) );
  NAND2X1 U8056 ( .A(ram[3876]), .B(n12793), .Y(n4198) );
  OAI21X1 U8057 ( .A(n12749), .B(n12793), .C(n4199), .Y(n8314) );
  NAND2X1 U8058 ( .A(ram[3877]), .B(n12793), .Y(n4199) );
  OAI21X1 U8059 ( .A(n12743), .B(n12793), .C(n4200), .Y(n8315) );
  NAND2X1 U8060 ( .A(ram[3878]), .B(n12793), .Y(n4200) );
  OAI21X1 U8061 ( .A(n12737), .B(n12793), .C(n4201), .Y(n8316) );
  NAND2X1 U8062 ( .A(ram[3879]), .B(n12793), .Y(n4201) );
  OAI21X1 U8063 ( .A(n12731), .B(n12793), .C(n4202), .Y(n8317) );
  NAND2X1 U8064 ( .A(ram[3880]), .B(n12793), .Y(n4202) );
  OAI21X1 U8065 ( .A(n12725), .B(n12793), .C(n4203), .Y(n8318) );
  NAND2X1 U8066 ( .A(ram[3881]), .B(n12793), .Y(n4203) );
  OAI21X1 U8067 ( .A(n12719), .B(n12793), .C(n4204), .Y(n8319) );
  NAND2X1 U8068 ( .A(ram[3882]), .B(n12793), .Y(n4204) );
  OAI21X1 U8069 ( .A(n12713), .B(n12793), .C(n4205), .Y(n8320) );
  NAND2X1 U8070 ( .A(ram[3883]), .B(n12793), .Y(n4205) );
  OAI21X1 U8071 ( .A(n12707), .B(n12793), .C(n4206), .Y(n8321) );
  NAND2X1 U8072 ( .A(ram[3884]), .B(n12793), .Y(n4206) );
  OAI21X1 U8073 ( .A(n12701), .B(n12793), .C(n4207), .Y(n8322) );
  NAND2X1 U8074 ( .A(ram[3885]), .B(n12793), .Y(n4207) );
  OAI21X1 U8075 ( .A(n12695), .B(n12793), .C(n4208), .Y(n8323) );
  NAND2X1 U8076 ( .A(ram[3886]), .B(n12793), .Y(n4208) );
  OAI21X1 U8077 ( .A(n12689), .B(n12793), .C(n4209), .Y(n8324) );
  NAND2X1 U8078 ( .A(ram[3887]), .B(n12793), .Y(n4209) );
  OAI21X1 U8081 ( .A(n12778), .B(n12792), .C(n4212), .Y(n8325) );
  NAND2X1 U8082 ( .A(ram[3888]), .B(n12792), .Y(n4212) );
  OAI21X1 U8083 ( .A(n12772), .B(n12792), .C(n4213), .Y(n8326) );
  NAND2X1 U8084 ( .A(ram[3889]), .B(n12792), .Y(n4213) );
  OAI21X1 U8085 ( .A(n12766), .B(n12792), .C(n4214), .Y(n8327) );
  NAND2X1 U8086 ( .A(ram[3890]), .B(n12792), .Y(n4214) );
  OAI21X1 U8087 ( .A(n12760), .B(n12792), .C(n4215), .Y(n8328) );
  NAND2X1 U8088 ( .A(ram[3891]), .B(n12792), .Y(n4215) );
  OAI21X1 U8089 ( .A(n12754), .B(n12792), .C(n4216), .Y(n8329) );
  NAND2X1 U8090 ( .A(ram[3892]), .B(n12792), .Y(n4216) );
  OAI21X1 U8091 ( .A(n12748), .B(n12792), .C(n4217), .Y(n8330) );
  NAND2X1 U8092 ( .A(ram[3893]), .B(n12792), .Y(n4217) );
  OAI21X1 U8093 ( .A(n12742), .B(n12792), .C(n4218), .Y(n8331) );
  NAND2X1 U8094 ( .A(ram[3894]), .B(n12792), .Y(n4218) );
  OAI21X1 U8095 ( .A(n12736), .B(n12792), .C(n4219), .Y(n8332) );
  NAND2X1 U8096 ( .A(ram[3895]), .B(n12792), .Y(n4219) );
  OAI21X1 U8097 ( .A(n12730), .B(n12792), .C(n4220), .Y(n8333) );
  NAND2X1 U8098 ( .A(ram[3896]), .B(n12792), .Y(n4220) );
  OAI21X1 U8099 ( .A(n12724), .B(n12792), .C(n4221), .Y(n8334) );
  NAND2X1 U8100 ( .A(ram[3897]), .B(n12792), .Y(n4221) );
  OAI21X1 U8101 ( .A(n12718), .B(n12792), .C(n4222), .Y(n8335) );
  NAND2X1 U8102 ( .A(ram[3898]), .B(n12792), .Y(n4222) );
  OAI21X1 U8103 ( .A(n12712), .B(n12792), .C(n4223), .Y(n8336) );
  NAND2X1 U8104 ( .A(ram[3899]), .B(n12792), .Y(n4223) );
  OAI21X1 U8105 ( .A(n12706), .B(n12792), .C(n4224), .Y(n8337) );
  NAND2X1 U8106 ( .A(ram[3900]), .B(n12792), .Y(n4224) );
  OAI21X1 U8107 ( .A(n12700), .B(n12792), .C(n4225), .Y(n8338) );
  NAND2X1 U8108 ( .A(ram[3901]), .B(n12792), .Y(n4225) );
  OAI21X1 U8109 ( .A(n12694), .B(n12792), .C(n4226), .Y(n8339) );
  NAND2X1 U8110 ( .A(ram[3902]), .B(n12792), .Y(n4226) );
  OAI21X1 U8111 ( .A(n12688), .B(n12792), .C(n4227), .Y(n8340) );
  NAND2X1 U8112 ( .A(ram[3903]), .B(n12792), .Y(n4227) );
  NOR2X1 U8115 ( .A(mem_access_addr[2]), .B(mem_access_addr[3]), .Y(n4173) );
  OAI21X1 U8116 ( .A(n12777), .B(n12791), .C(n4230), .Y(n8341) );
  NAND2X1 U8117 ( .A(ram[3904]), .B(n12791), .Y(n4230) );
  OAI21X1 U8118 ( .A(n12771), .B(n12791), .C(n4231), .Y(n8342) );
  NAND2X1 U8119 ( .A(ram[3905]), .B(n12791), .Y(n4231) );
  OAI21X1 U8120 ( .A(n12765), .B(n12791), .C(n4232), .Y(n8343) );
  NAND2X1 U8121 ( .A(ram[3906]), .B(n12791), .Y(n4232) );
  OAI21X1 U8122 ( .A(n12759), .B(n12791), .C(n4233), .Y(n8344) );
  NAND2X1 U8123 ( .A(ram[3907]), .B(n12791), .Y(n4233) );
  OAI21X1 U8124 ( .A(n12753), .B(n12791), .C(n4234), .Y(n8345) );
  NAND2X1 U8125 ( .A(ram[3908]), .B(n12791), .Y(n4234) );
  OAI21X1 U8126 ( .A(n12747), .B(n12791), .C(n4235), .Y(n8346) );
  NAND2X1 U8127 ( .A(ram[3909]), .B(n12791), .Y(n4235) );
  OAI21X1 U8128 ( .A(n12741), .B(n12791), .C(n4236), .Y(n8347) );
  NAND2X1 U8129 ( .A(ram[3910]), .B(n12791), .Y(n4236) );
  OAI21X1 U8130 ( .A(n12735), .B(n12791), .C(n4237), .Y(n8348) );
  NAND2X1 U8131 ( .A(ram[3911]), .B(n12791), .Y(n4237) );
  OAI21X1 U8132 ( .A(n12729), .B(n12791), .C(n4238), .Y(n8349) );
  NAND2X1 U8133 ( .A(ram[3912]), .B(n12791), .Y(n4238) );
  OAI21X1 U8134 ( .A(n12723), .B(n12791), .C(n4239), .Y(n8350) );
  NAND2X1 U8135 ( .A(ram[3913]), .B(n12791), .Y(n4239) );
  OAI21X1 U8136 ( .A(n12717), .B(n12791), .C(n4240), .Y(n8351) );
  NAND2X1 U8137 ( .A(ram[3914]), .B(n12791), .Y(n4240) );
  OAI21X1 U8138 ( .A(n12711), .B(n12791), .C(n4241), .Y(n8352) );
  NAND2X1 U8139 ( .A(ram[3915]), .B(n12791), .Y(n4241) );
  OAI21X1 U8140 ( .A(n12705), .B(n12791), .C(n4242), .Y(n8353) );
  NAND2X1 U8141 ( .A(ram[3916]), .B(n12791), .Y(n4242) );
  OAI21X1 U8142 ( .A(n12699), .B(n12791), .C(n4243), .Y(n8354) );
  NAND2X1 U8143 ( .A(ram[3917]), .B(n12791), .Y(n4243) );
  OAI21X1 U8144 ( .A(n12693), .B(n12791), .C(n4244), .Y(n8355) );
  NAND2X1 U8145 ( .A(ram[3918]), .B(n12791), .Y(n4244) );
  OAI21X1 U8146 ( .A(n12687), .B(n12791), .C(n4245), .Y(n8356) );
  NAND2X1 U8147 ( .A(ram[3919]), .B(n12791), .Y(n4245) );
  OAI21X1 U8150 ( .A(n12776), .B(n12790), .C(n4248), .Y(n8357) );
  NAND2X1 U8151 ( .A(ram[3920]), .B(n12790), .Y(n4248) );
  OAI21X1 U8152 ( .A(n12770), .B(n12790), .C(n4249), .Y(n8358) );
  NAND2X1 U8153 ( .A(ram[3921]), .B(n12790), .Y(n4249) );
  OAI21X1 U8154 ( .A(n12764), .B(n12790), .C(n4250), .Y(n8359) );
  NAND2X1 U8155 ( .A(ram[3922]), .B(n12790), .Y(n4250) );
  OAI21X1 U8156 ( .A(n12758), .B(n12790), .C(n4251), .Y(n8360) );
  NAND2X1 U8157 ( .A(ram[3923]), .B(n12790), .Y(n4251) );
  OAI21X1 U8158 ( .A(n12752), .B(n12790), .C(n4252), .Y(n8361) );
  NAND2X1 U8159 ( .A(ram[3924]), .B(n12790), .Y(n4252) );
  OAI21X1 U8160 ( .A(n12746), .B(n12790), .C(n4253), .Y(n8362) );
  NAND2X1 U8161 ( .A(ram[3925]), .B(n12790), .Y(n4253) );
  OAI21X1 U8162 ( .A(n12740), .B(n12790), .C(n4254), .Y(n8363) );
  NAND2X1 U8163 ( .A(ram[3926]), .B(n12790), .Y(n4254) );
  OAI21X1 U8164 ( .A(n12734), .B(n12790), .C(n4255), .Y(n8364) );
  NAND2X1 U8165 ( .A(ram[3927]), .B(n12790), .Y(n4255) );
  OAI21X1 U8166 ( .A(n12728), .B(n12790), .C(n4256), .Y(n8365) );
  NAND2X1 U8167 ( .A(ram[3928]), .B(n12790), .Y(n4256) );
  OAI21X1 U8168 ( .A(n12722), .B(n12790), .C(n4257), .Y(n8366) );
  NAND2X1 U8169 ( .A(ram[3929]), .B(n12790), .Y(n4257) );
  OAI21X1 U8170 ( .A(n12716), .B(n12790), .C(n4258), .Y(n8367) );
  NAND2X1 U8171 ( .A(ram[3930]), .B(n12790), .Y(n4258) );
  OAI21X1 U8172 ( .A(n12710), .B(n12790), .C(n4259), .Y(n8368) );
  NAND2X1 U8173 ( .A(ram[3931]), .B(n12790), .Y(n4259) );
  OAI21X1 U8174 ( .A(n12704), .B(n12790), .C(n4260), .Y(n8369) );
  NAND2X1 U8175 ( .A(ram[3932]), .B(n12790), .Y(n4260) );
  OAI21X1 U8176 ( .A(n12698), .B(n12790), .C(n4261), .Y(n8370) );
  NAND2X1 U8177 ( .A(ram[3933]), .B(n12790), .Y(n4261) );
  OAI21X1 U8178 ( .A(n12692), .B(n12790), .C(n4262), .Y(n8371) );
  NAND2X1 U8179 ( .A(ram[3934]), .B(n12790), .Y(n4262) );
  OAI21X1 U8180 ( .A(n12686), .B(n12790), .C(n4263), .Y(n8372) );
  NAND2X1 U8181 ( .A(ram[3935]), .B(n12790), .Y(n4263) );
  OAI21X1 U8184 ( .A(n12779), .B(n12789), .C(n4265), .Y(n8373) );
  NAND2X1 U8185 ( .A(ram[3936]), .B(n12789), .Y(n4265) );
  OAI21X1 U8186 ( .A(n12773), .B(n12789), .C(n4266), .Y(n8374) );
  NAND2X1 U8187 ( .A(ram[3937]), .B(n12789), .Y(n4266) );
  OAI21X1 U8188 ( .A(n12767), .B(n12789), .C(n4267), .Y(n8375) );
  NAND2X1 U8189 ( .A(ram[3938]), .B(n12789), .Y(n4267) );
  OAI21X1 U8190 ( .A(n12761), .B(n12789), .C(n4268), .Y(n8376) );
  NAND2X1 U8191 ( .A(ram[3939]), .B(n12789), .Y(n4268) );
  OAI21X1 U8192 ( .A(n12755), .B(n12789), .C(n4269), .Y(n8377) );
  NAND2X1 U8193 ( .A(ram[3940]), .B(n12789), .Y(n4269) );
  OAI21X1 U8194 ( .A(n12749), .B(n12789), .C(n4270), .Y(n8378) );
  NAND2X1 U8195 ( .A(ram[3941]), .B(n12789), .Y(n4270) );
  OAI21X1 U8196 ( .A(n12743), .B(n12789), .C(n4271), .Y(n8379) );
  NAND2X1 U8197 ( .A(ram[3942]), .B(n12789), .Y(n4271) );
  OAI21X1 U8198 ( .A(n12737), .B(n12789), .C(n4272), .Y(n8380) );
  NAND2X1 U8199 ( .A(ram[3943]), .B(n12789), .Y(n4272) );
  OAI21X1 U8200 ( .A(n12731), .B(n12789), .C(n4273), .Y(n8381) );
  NAND2X1 U8201 ( .A(ram[3944]), .B(n12789), .Y(n4273) );
  OAI21X1 U8202 ( .A(n12725), .B(n12789), .C(n4274), .Y(n8382) );
  NAND2X1 U8203 ( .A(ram[3945]), .B(n12789), .Y(n4274) );
  OAI21X1 U8204 ( .A(n12719), .B(n12789), .C(n4275), .Y(n8383) );
  NAND2X1 U8205 ( .A(ram[3946]), .B(n12789), .Y(n4275) );
  OAI21X1 U8206 ( .A(n12713), .B(n12789), .C(n4276), .Y(n8384) );
  NAND2X1 U8207 ( .A(ram[3947]), .B(n12789), .Y(n4276) );
  OAI21X1 U8208 ( .A(n12707), .B(n12789), .C(n4277), .Y(n8385) );
  NAND2X1 U8209 ( .A(ram[3948]), .B(n12789), .Y(n4277) );
  OAI21X1 U8210 ( .A(n12701), .B(n12789), .C(n4278), .Y(n8386) );
  NAND2X1 U8211 ( .A(ram[3949]), .B(n12789), .Y(n4278) );
  OAI21X1 U8212 ( .A(n12695), .B(n12789), .C(n4279), .Y(n8387) );
  NAND2X1 U8213 ( .A(ram[3950]), .B(n12789), .Y(n4279) );
  OAI21X1 U8214 ( .A(n12689), .B(n12789), .C(n4280), .Y(n8388) );
  NAND2X1 U8215 ( .A(ram[3951]), .B(n12789), .Y(n4280) );
  OAI21X1 U8218 ( .A(n12777), .B(n12788), .C(n4282), .Y(n8389) );
  NAND2X1 U8219 ( .A(ram[3952]), .B(n12788), .Y(n4282) );
  OAI21X1 U8220 ( .A(n12771), .B(n12788), .C(n4283), .Y(n8390) );
  NAND2X1 U8221 ( .A(ram[3953]), .B(n12788), .Y(n4283) );
  OAI21X1 U8222 ( .A(n12764), .B(n12788), .C(n4284), .Y(n8391) );
  NAND2X1 U8223 ( .A(ram[3954]), .B(n12788), .Y(n4284) );
  OAI21X1 U8224 ( .A(n12758), .B(n12788), .C(n4285), .Y(n8392) );
  NAND2X1 U8225 ( .A(ram[3955]), .B(n12788), .Y(n4285) );
  OAI21X1 U8226 ( .A(n12752), .B(n12788), .C(n4286), .Y(n8393) );
  NAND2X1 U8227 ( .A(ram[3956]), .B(n12788), .Y(n4286) );
  OAI21X1 U8228 ( .A(n12746), .B(n12788), .C(n4287), .Y(n8394) );
  NAND2X1 U8229 ( .A(ram[3957]), .B(n12788), .Y(n4287) );
  OAI21X1 U8230 ( .A(n12740), .B(n12788), .C(n4288), .Y(n8395) );
  NAND2X1 U8231 ( .A(ram[3958]), .B(n12788), .Y(n4288) );
  OAI21X1 U8232 ( .A(n12734), .B(n12788), .C(n4289), .Y(n8396) );
  NAND2X1 U8233 ( .A(ram[3959]), .B(n12788), .Y(n4289) );
  OAI21X1 U8234 ( .A(n12728), .B(n12788), .C(n4290), .Y(n8397) );
  NAND2X1 U8235 ( .A(ram[3960]), .B(n12788), .Y(n4290) );
  OAI21X1 U8236 ( .A(n12722), .B(n12788), .C(n4291), .Y(n8398) );
  NAND2X1 U8237 ( .A(ram[3961]), .B(n12788), .Y(n4291) );
  OAI21X1 U8238 ( .A(n12716), .B(n12788), .C(n4292), .Y(n8399) );
  NAND2X1 U8239 ( .A(ram[3962]), .B(n12788), .Y(n4292) );
  OAI21X1 U8240 ( .A(n12710), .B(n12788), .C(n4293), .Y(n8400) );
  NAND2X1 U8241 ( .A(ram[3963]), .B(n12788), .Y(n4293) );
  OAI21X1 U8242 ( .A(n12704), .B(n12788), .C(n4294), .Y(n8401) );
  NAND2X1 U8243 ( .A(ram[3964]), .B(n12788), .Y(n4294) );
  OAI21X1 U8244 ( .A(n12698), .B(n12788), .C(n4295), .Y(n8402) );
  NAND2X1 U8245 ( .A(ram[3965]), .B(n12788), .Y(n4295) );
  OAI21X1 U8246 ( .A(n12693), .B(n12788), .C(n4296), .Y(n8403) );
  NAND2X1 U8247 ( .A(ram[3966]), .B(n12788), .Y(n4296) );
  OAI21X1 U8248 ( .A(n12687), .B(n12788), .C(n4297), .Y(n8404) );
  NAND2X1 U8249 ( .A(ram[3967]), .B(n12788), .Y(n4297) );
  NOR2X1 U8252 ( .A(n13037), .B(mem_access_addr[3]), .Y(n4246) );
  OAI21X1 U8253 ( .A(n12776), .B(n12787), .C(n4299), .Y(n8405) );
  NAND2X1 U8254 ( .A(ram[3968]), .B(n12787), .Y(n4299) );
  OAI21X1 U8255 ( .A(n12770), .B(n12787), .C(n4300), .Y(n8406) );
  NAND2X1 U8256 ( .A(ram[3969]), .B(n12787), .Y(n4300) );
  OAI21X1 U8257 ( .A(n12765), .B(n12787), .C(n4301), .Y(n8407) );
  NAND2X1 U8258 ( .A(ram[3970]), .B(n12787), .Y(n4301) );
  OAI21X1 U8259 ( .A(n12759), .B(n12787), .C(n4302), .Y(n8408) );
  NAND2X1 U8260 ( .A(ram[3971]), .B(n12787), .Y(n4302) );
  OAI21X1 U8261 ( .A(n12753), .B(n12787), .C(n4303), .Y(n8409) );
  NAND2X1 U8262 ( .A(ram[3972]), .B(n12787), .Y(n4303) );
  OAI21X1 U8263 ( .A(n12747), .B(n12787), .C(n4304), .Y(n8410) );
  NAND2X1 U8264 ( .A(ram[3973]), .B(n12787), .Y(n4304) );
  OAI21X1 U8265 ( .A(n12741), .B(n12787), .C(n4305), .Y(n8411) );
  NAND2X1 U8266 ( .A(ram[3974]), .B(n12787), .Y(n4305) );
  OAI21X1 U8267 ( .A(n12735), .B(n12787), .C(n4306), .Y(n8412) );
  NAND2X1 U8268 ( .A(ram[3975]), .B(n12787), .Y(n4306) );
  OAI21X1 U8269 ( .A(n12729), .B(n12787), .C(n4307), .Y(n8413) );
  NAND2X1 U8270 ( .A(ram[3976]), .B(n12787), .Y(n4307) );
  OAI21X1 U8271 ( .A(n12723), .B(n12787), .C(n4308), .Y(n8414) );
  NAND2X1 U8272 ( .A(ram[3977]), .B(n12787), .Y(n4308) );
  OAI21X1 U8273 ( .A(n12717), .B(n12787), .C(n4309), .Y(n8415) );
  NAND2X1 U8274 ( .A(ram[3978]), .B(n12787), .Y(n4309) );
  OAI21X1 U8275 ( .A(n12711), .B(n12787), .C(n4310), .Y(n8416) );
  NAND2X1 U8276 ( .A(ram[3979]), .B(n12787), .Y(n4310) );
  OAI21X1 U8277 ( .A(n12705), .B(n12787), .C(n4311), .Y(n8417) );
  NAND2X1 U8278 ( .A(ram[3980]), .B(n12787), .Y(n4311) );
  OAI21X1 U8279 ( .A(n12699), .B(n12787), .C(n4312), .Y(n8418) );
  NAND2X1 U8280 ( .A(ram[3981]), .B(n12787), .Y(n4312) );
  OAI21X1 U8281 ( .A(n12692), .B(n12787), .C(n4313), .Y(n8419) );
  NAND2X1 U8282 ( .A(ram[3982]), .B(n12787), .Y(n4313) );
  OAI21X1 U8283 ( .A(n12686), .B(n12787), .C(n4314), .Y(n8420) );
  NAND2X1 U8284 ( .A(ram[3983]), .B(n12787), .Y(n4314) );
  OAI21X1 U8287 ( .A(n12777), .B(n12786), .C(n4317), .Y(n8421) );
  NAND2X1 U8288 ( .A(ram[3984]), .B(n12786), .Y(n4317) );
  OAI21X1 U8289 ( .A(n12771), .B(n12786), .C(n4318), .Y(n8422) );
  NAND2X1 U8290 ( .A(ram[3985]), .B(n12786), .Y(n4318) );
  OAI21X1 U8291 ( .A(n12766), .B(n12786), .C(n4319), .Y(n8423) );
  NAND2X1 U8292 ( .A(ram[3986]), .B(n12786), .Y(n4319) );
  OAI21X1 U8293 ( .A(n12760), .B(n12786), .C(n4320), .Y(n8424) );
  NAND2X1 U8294 ( .A(ram[3987]), .B(n12786), .Y(n4320) );
  OAI21X1 U8295 ( .A(n12754), .B(n12786), .C(n4321), .Y(n8425) );
  NAND2X1 U8296 ( .A(ram[3988]), .B(n12786), .Y(n4321) );
  OAI21X1 U8297 ( .A(n12748), .B(n12786), .C(n4322), .Y(n8426) );
  NAND2X1 U8298 ( .A(ram[3989]), .B(n12786), .Y(n4322) );
  OAI21X1 U8299 ( .A(n12742), .B(n12786), .C(n4323), .Y(n8427) );
  NAND2X1 U8300 ( .A(ram[3990]), .B(n12786), .Y(n4323) );
  OAI21X1 U8301 ( .A(n12736), .B(n12786), .C(n4324), .Y(n8428) );
  NAND2X1 U8302 ( .A(ram[3991]), .B(n12786), .Y(n4324) );
  OAI21X1 U8303 ( .A(n12730), .B(n12786), .C(n4325), .Y(n8429) );
  NAND2X1 U8304 ( .A(ram[3992]), .B(n12786), .Y(n4325) );
  OAI21X1 U8305 ( .A(n12724), .B(n12786), .C(n4326), .Y(n8430) );
  NAND2X1 U8306 ( .A(ram[3993]), .B(n12786), .Y(n4326) );
  OAI21X1 U8307 ( .A(n12718), .B(n12786), .C(n4327), .Y(n8431) );
  NAND2X1 U8308 ( .A(ram[3994]), .B(n12786), .Y(n4327) );
  OAI21X1 U8309 ( .A(n12712), .B(n12786), .C(n4328), .Y(n8432) );
  NAND2X1 U8310 ( .A(ram[3995]), .B(n12786), .Y(n4328) );
  OAI21X1 U8311 ( .A(n12706), .B(n12786), .C(n4329), .Y(n8433) );
  NAND2X1 U8312 ( .A(ram[3996]), .B(n12786), .Y(n4329) );
  OAI21X1 U8313 ( .A(n12700), .B(n12786), .C(n4330), .Y(n8434) );
  NAND2X1 U8314 ( .A(ram[3997]), .B(n12786), .Y(n4330) );
  OAI21X1 U8315 ( .A(n12693), .B(n12786), .C(n4331), .Y(n8435) );
  NAND2X1 U8316 ( .A(ram[3998]), .B(n12786), .Y(n4331) );
  OAI21X1 U8317 ( .A(n12687), .B(n12786), .C(n4332), .Y(n8436) );
  NAND2X1 U8318 ( .A(ram[3999]), .B(n12786), .Y(n4332) );
  OAI21X1 U8321 ( .A(n12779), .B(n12785), .C(n4334), .Y(n8437) );
  NAND2X1 U8322 ( .A(ram[4000]), .B(n12785), .Y(n4334) );
  OAI21X1 U8323 ( .A(n12773), .B(n12785), .C(n4335), .Y(n8438) );
  NAND2X1 U8324 ( .A(ram[4001]), .B(n12785), .Y(n4335) );
  OAI21X1 U8325 ( .A(n12765), .B(n12785), .C(n4336), .Y(n8439) );
  NAND2X1 U8326 ( .A(ram[4002]), .B(n12785), .Y(n4336) );
  OAI21X1 U8327 ( .A(n12759), .B(n12785), .C(n4337), .Y(n8440) );
  NAND2X1 U8328 ( .A(ram[4003]), .B(n12785), .Y(n4337) );
  OAI21X1 U8329 ( .A(n12753), .B(n12785), .C(n4338), .Y(n8441) );
  NAND2X1 U8330 ( .A(ram[4004]), .B(n12785), .Y(n4338) );
  OAI21X1 U8331 ( .A(n12747), .B(n12785), .C(n4339), .Y(n8442) );
  NAND2X1 U8332 ( .A(ram[4005]), .B(n12785), .Y(n4339) );
  OAI21X1 U8333 ( .A(n12741), .B(n12785), .C(n4340), .Y(n8443) );
  NAND2X1 U8334 ( .A(ram[4006]), .B(n12785), .Y(n4340) );
  OAI21X1 U8335 ( .A(n12735), .B(n12785), .C(n4341), .Y(n8444) );
  NAND2X1 U8336 ( .A(ram[4007]), .B(n12785), .Y(n4341) );
  OAI21X1 U8337 ( .A(n12729), .B(n12785), .C(n4342), .Y(n8445) );
  NAND2X1 U8338 ( .A(ram[4008]), .B(n12785), .Y(n4342) );
  OAI21X1 U8339 ( .A(n12723), .B(n12785), .C(n4343), .Y(n8446) );
  NAND2X1 U8340 ( .A(ram[4009]), .B(n12785), .Y(n4343) );
  OAI21X1 U8341 ( .A(n12717), .B(n12785), .C(n4344), .Y(n8447) );
  NAND2X1 U8342 ( .A(ram[4010]), .B(n12785), .Y(n4344) );
  OAI21X1 U8343 ( .A(n12711), .B(n12785), .C(n4345), .Y(n8448) );
  NAND2X1 U8344 ( .A(ram[4011]), .B(n12785), .Y(n4345) );
  OAI21X1 U8345 ( .A(n12705), .B(n12785), .C(n4346), .Y(n8449) );
  NAND2X1 U8346 ( .A(ram[4012]), .B(n12785), .Y(n4346) );
  OAI21X1 U8347 ( .A(n12699), .B(n12785), .C(n4347), .Y(n8450) );
  NAND2X1 U8348 ( .A(ram[4013]), .B(n12785), .Y(n4347) );
  OAI21X1 U8349 ( .A(n12695), .B(n12785), .C(n4348), .Y(n8451) );
  NAND2X1 U8350 ( .A(ram[4014]), .B(n12785), .Y(n4348) );
  OAI21X1 U8351 ( .A(n12689), .B(n12785), .C(n4349), .Y(n8452) );
  NAND2X1 U8352 ( .A(ram[4015]), .B(n12785), .Y(n4349) );
  OAI21X1 U8355 ( .A(n12778), .B(n12784), .C(n4351), .Y(n8453) );
  NAND2X1 U8356 ( .A(ram[4016]), .B(n12784), .Y(n4351) );
  OAI21X1 U8357 ( .A(n12772), .B(n12784), .C(n4352), .Y(n8454) );
  NAND2X1 U8358 ( .A(ram[4017]), .B(n12784), .Y(n4352) );
  OAI21X1 U8359 ( .A(n12767), .B(n12784), .C(n4353), .Y(n8455) );
  NAND2X1 U8360 ( .A(ram[4018]), .B(n12784), .Y(n4353) );
  OAI21X1 U8361 ( .A(n12761), .B(n12784), .C(n4354), .Y(n8456) );
  NAND2X1 U8362 ( .A(ram[4019]), .B(n12784), .Y(n4354) );
  OAI21X1 U8363 ( .A(n12755), .B(n12784), .C(n4355), .Y(n8457) );
  NAND2X1 U8364 ( .A(ram[4020]), .B(n12784), .Y(n4355) );
  OAI21X1 U8365 ( .A(n12749), .B(n12784), .C(n4356), .Y(n8458) );
  NAND2X1 U8366 ( .A(ram[4021]), .B(n12784), .Y(n4356) );
  OAI21X1 U8367 ( .A(n12743), .B(n12784), .C(n4357), .Y(n8459) );
  NAND2X1 U8368 ( .A(ram[4022]), .B(n12784), .Y(n4357) );
  OAI21X1 U8369 ( .A(n12737), .B(n12784), .C(n4358), .Y(n8460) );
  NAND2X1 U8370 ( .A(ram[4023]), .B(n12784), .Y(n4358) );
  OAI21X1 U8371 ( .A(n12731), .B(n12784), .C(n4359), .Y(n8461) );
  NAND2X1 U8372 ( .A(ram[4024]), .B(n12784), .Y(n4359) );
  OAI21X1 U8373 ( .A(n12725), .B(n12784), .C(n4360), .Y(n8462) );
  NAND2X1 U8374 ( .A(ram[4025]), .B(n12784), .Y(n4360) );
  OAI21X1 U8375 ( .A(n12719), .B(n12784), .C(n4361), .Y(n8463) );
  NAND2X1 U8376 ( .A(ram[4026]), .B(n12784), .Y(n4361) );
  OAI21X1 U8377 ( .A(n12713), .B(n12784), .C(n4362), .Y(n8464) );
  NAND2X1 U8378 ( .A(ram[4027]), .B(n12784), .Y(n4362) );
  OAI21X1 U8379 ( .A(n12707), .B(n12784), .C(n4363), .Y(n8465) );
  NAND2X1 U8380 ( .A(ram[4028]), .B(n12784), .Y(n4363) );
  OAI21X1 U8381 ( .A(n12701), .B(n12784), .C(n4364), .Y(n8466) );
  NAND2X1 U8382 ( .A(ram[4029]), .B(n12784), .Y(n4364) );
  OAI21X1 U8383 ( .A(n12694), .B(n12784), .C(n4365), .Y(n8467) );
  NAND2X1 U8384 ( .A(ram[4030]), .B(n12784), .Y(n4365) );
  OAI21X1 U8385 ( .A(n12688), .B(n12784), .C(n4366), .Y(n8468) );
  NAND2X1 U8386 ( .A(ram[4031]), .B(n12784), .Y(n4366) );
  AND2X1 U8389 ( .A(mem_access_addr[3]), .B(n13037), .Y(n4315) );
  OAI21X1 U8390 ( .A(n12776), .B(n12783), .C(n4368), .Y(n8469) );
  NAND2X1 U8391 ( .A(ram[4032]), .B(n12783), .Y(n4368) );
  OAI21X1 U8392 ( .A(n12770), .B(n12783), .C(n4369), .Y(n8470) );
  NAND2X1 U8393 ( .A(ram[4033]), .B(n12783), .Y(n4369) );
  OAI21X1 U8394 ( .A(n12764), .B(n12783), .C(n4370), .Y(n8471) );
  NAND2X1 U8395 ( .A(ram[4034]), .B(n12783), .Y(n4370) );
  OAI21X1 U8396 ( .A(n12758), .B(n12783), .C(n4371), .Y(n8472) );
  NAND2X1 U8397 ( .A(ram[4035]), .B(n12783), .Y(n4371) );
  OAI21X1 U8398 ( .A(n12752), .B(n12783), .C(n4372), .Y(n8473) );
  NAND2X1 U8399 ( .A(ram[4036]), .B(n12783), .Y(n4372) );
  OAI21X1 U8400 ( .A(n12746), .B(n12783), .C(n4373), .Y(n8474) );
  NAND2X1 U8401 ( .A(ram[4037]), .B(n12783), .Y(n4373) );
  OAI21X1 U8402 ( .A(n12740), .B(n12783), .C(n4374), .Y(n8475) );
  NAND2X1 U8403 ( .A(ram[4038]), .B(n12783), .Y(n4374) );
  OAI21X1 U8404 ( .A(n12734), .B(n12783), .C(n4375), .Y(n8476) );
  NAND2X1 U8405 ( .A(ram[4039]), .B(n12783), .Y(n4375) );
  OAI21X1 U8406 ( .A(n12728), .B(n12783), .C(n4376), .Y(n8477) );
  NAND2X1 U8407 ( .A(ram[4040]), .B(n12783), .Y(n4376) );
  OAI21X1 U8408 ( .A(n12722), .B(n12783), .C(n4377), .Y(n8478) );
  NAND2X1 U8409 ( .A(ram[4041]), .B(n12783), .Y(n4377) );
  OAI21X1 U8410 ( .A(n12716), .B(n12783), .C(n4378), .Y(n8479) );
  NAND2X1 U8411 ( .A(ram[4042]), .B(n12783), .Y(n4378) );
  OAI21X1 U8412 ( .A(n12710), .B(n12783), .C(n4379), .Y(n8480) );
  NAND2X1 U8413 ( .A(ram[4043]), .B(n12783), .Y(n4379) );
  OAI21X1 U8414 ( .A(n12704), .B(n12783), .C(n4380), .Y(n8481) );
  NAND2X1 U8415 ( .A(ram[4044]), .B(n12783), .Y(n4380) );
  OAI21X1 U8416 ( .A(n12698), .B(n12783), .C(n4381), .Y(n8482) );
  NAND2X1 U8417 ( .A(ram[4045]), .B(n12783), .Y(n4381) );
  OAI21X1 U8418 ( .A(n12692), .B(n12783), .C(n4382), .Y(n8483) );
  NAND2X1 U8419 ( .A(ram[4046]), .B(n12783), .Y(n4382) );
  OAI21X1 U8420 ( .A(n12686), .B(n12783), .C(n4383), .Y(n8484) );
  NAND2X1 U8421 ( .A(ram[4047]), .B(n12783), .Y(n4383) );
  NOR2X1 U8424 ( .A(mem_access_addr[0]), .B(mem_access_addr[1]), .Y(n4174) );
  OAI21X1 U8425 ( .A(n12776), .B(n12782), .C(n4386), .Y(n8485) );
  NAND2X1 U8426 ( .A(ram[4048]), .B(n12782), .Y(n4386) );
  OAI21X1 U8427 ( .A(n12770), .B(n12782), .C(n4387), .Y(n8486) );
  NAND2X1 U8428 ( .A(ram[4049]), .B(n12782), .Y(n4387) );
  OAI21X1 U8429 ( .A(n12764), .B(n12782), .C(n4388), .Y(n8487) );
  NAND2X1 U8430 ( .A(ram[4050]), .B(n12782), .Y(n4388) );
  OAI21X1 U8431 ( .A(n12758), .B(n12782), .C(n4389), .Y(n8488) );
  NAND2X1 U8432 ( .A(ram[4051]), .B(n12782), .Y(n4389) );
  OAI21X1 U8433 ( .A(n12752), .B(n12782), .C(n4390), .Y(n8489) );
  NAND2X1 U8434 ( .A(ram[4052]), .B(n12782), .Y(n4390) );
  OAI21X1 U8435 ( .A(n12746), .B(n12782), .C(n4391), .Y(n8490) );
  NAND2X1 U8436 ( .A(ram[4053]), .B(n12782), .Y(n4391) );
  OAI21X1 U8437 ( .A(n12740), .B(n12782), .C(n4392), .Y(n8491) );
  NAND2X1 U8438 ( .A(ram[4054]), .B(n12782), .Y(n4392) );
  OAI21X1 U8439 ( .A(n12734), .B(n12782), .C(n4393), .Y(n8492) );
  NAND2X1 U8440 ( .A(ram[4055]), .B(n12782), .Y(n4393) );
  OAI21X1 U8441 ( .A(n12728), .B(n12782), .C(n4394), .Y(n8493) );
  NAND2X1 U8442 ( .A(ram[4056]), .B(n12782), .Y(n4394) );
  OAI21X1 U8443 ( .A(n12722), .B(n12782), .C(n4395), .Y(n8494) );
  NAND2X1 U8444 ( .A(ram[4057]), .B(n12782), .Y(n4395) );
  OAI21X1 U8445 ( .A(n12716), .B(n12782), .C(n4396), .Y(n8495) );
  NAND2X1 U8446 ( .A(ram[4058]), .B(n12782), .Y(n4396) );
  OAI21X1 U8447 ( .A(n12710), .B(n12782), .C(n4397), .Y(n8496) );
  NAND2X1 U8448 ( .A(ram[4059]), .B(n12782), .Y(n4397) );
  OAI21X1 U8449 ( .A(n12704), .B(n12782), .C(n4398), .Y(n8497) );
  NAND2X1 U8450 ( .A(ram[4060]), .B(n12782), .Y(n4398) );
  OAI21X1 U8451 ( .A(n12698), .B(n12782), .C(n4399), .Y(n8498) );
  NAND2X1 U8452 ( .A(ram[4061]), .B(n12782), .Y(n4399) );
  OAI21X1 U8453 ( .A(n12692), .B(n12782), .C(n4400), .Y(n8499) );
  NAND2X1 U8454 ( .A(ram[4062]), .B(n12782), .Y(n4400) );
  OAI21X1 U8455 ( .A(n12686), .B(n12782), .C(n4401), .Y(n8500) );
  NAND2X1 U8456 ( .A(ram[4063]), .B(n12782), .Y(n4401) );
  NOR2X1 U8459 ( .A(n13036), .B(mem_access_addr[1]), .Y(n4192) );
  OAI21X1 U8460 ( .A(n12777), .B(n12781), .C(n4403), .Y(n8501) );
  NAND2X1 U8461 ( .A(ram[4064]), .B(n12781), .Y(n4403) );
  OAI21X1 U8462 ( .A(n12771), .B(n12781), .C(n4404), .Y(n8502) );
  NAND2X1 U8463 ( .A(ram[4065]), .B(n12781), .Y(n4404) );
  OAI21X1 U8464 ( .A(n12766), .B(n12781), .C(n4405), .Y(n8503) );
  NAND2X1 U8465 ( .A(ram[4066]), .B(n12781), .Y(n4405) );
  OAI21X1 U8466 ( .A(n12760), .B(n12781), .C(n4406), .Y(n8504) );
  NAND2X1 U8467 ( .A(ram[4067]), .B(n12781), .Y(n4406) );
  OAI21X1 U8468 ( .A(n12754), .B(n12781), .C(n4407), .Y(n8505) );
  NAND2X1 U8469 ( .A(ram[4068]), .B(n12781), .Y(n4407) );
  OAI21X1 U8470 ( .A(n12748), .B(n12781), .C(n4408), .Y(n8506) );
  NAND2X1 U8471 ( .A(ram[4069]), .B(n12781), .Y(n4408) );
  OAI21X1 U8472 ( .A(n12742), .B(n12781), .C(n4409), .Y(n8507) );
  NAND2X1 U8473 ( .A(ram[4070]), .B(n12781), .Y(n4409) );
  OAI21X1 U8474 ( .A(n12736), .B(n12781), .C(n4410), .Y(n8508) );
  NAND2X1 U8475 ( .A(ram[4071]), .B(n12781), .Y(n4410) );
  OAI21X1 U8476 ( .A(n12730), .B(n12781), .C(n4411), .Y(n8509) );
  NAND2X1 U8477 ( .A(ram[4072]), .B(n12781), .Y(n4411) );
  OAI21X1 U8478 ( .A(n12724), .B(n12781), .C(n4412), .Y(n8510) );
  NAND2X1 U8479 ( .A(ram[4073]), .B(n12781), .Y(n4412) );
  OAI21X1 U8480 ( .A(n12718), .B(n12781), .C(n4413), .Y(n8511) );
  NAND2X1 U8481 ( .A(ram[4074]), .B(n12781), .Y(n4413) );
  OAI21X1 U8482 ( .A(n12712), .B(n12781), .C(n4414), .Y(n8512) );
  NAND2X1 U8483 ( .A(ram[4075]), .B(n12781), .Y(n4414) );
  OAI21X1 U8484 ( .A(n12706), .B(n12781), .C(n4415), .Y(n8513) );
  NAND2X1 U8485 ( .A(ram[4076]), .B(n12781), .Y(n4415) );
  OAI21X1 U8486 ( .A(n12700), .B(n12781), .C(n4416), .Y(n8514) );
  NAND2X1 U8487 ( .A(ram[4077]), .B(n12781), .Y(n4416) );
  OAI21X1 U8488 ( .A(n12693), .B(n12781), .C(n4417), .Y(n8515) );
  NAND2X1 U8489 ( .A(ram[4078]), .B(n12781), .Y(n4417) );
  OAI21X1 U8490 ( .A(n12687), .B(n12781), .C(n4418), .Y(n8516) );
  NAND2X1 U8491 ( .A(ram[4079]), .B(n12781), .Y(n4418) );
  AND2X1 U8494 ( .A(mem_access_addr[1]), .B(n13036), .Y(n4210) );
  OAI21X1 U8495 ( .A(n12779), .B(n12780), .C(n4420), .Y(n8517) );
  NAND2X1 U8496 ( .A(ram[4080]), .B(n12780), .Y(n4420) );
  OAI21X1 U8497 ( .A(n12773), .B(n12780), .C(n4421), .Y(n8518) );
  NAND2X1 U8498 ( .A(ram[4081]), .B(n12780), .Y(n4421) );
  OAI21X1 U8499 ( .A(n12765), .B(n12780), .C(n4422), .Y(n8519) );
  NAND2X1 U8500 ( .A(ram[4082]), .B(n12780), .Y(n4422) );
  OAI21X1 U8501 ( .A(n12759), .B(n12780), .C(n4423), .Y(n8520) );
  NAND2X1 U8502 ( .A(ram[4083]), .B(n12780), .Y(n4423) );
  OAI21X1 U8503 ( .A(n12753), .B(n12780), .C(n4424), .Y(n8521) );
  NAND2X1 U8504 ( .A(ram[4084]), .B(n12780), .Y(n4424) );
  OAI21X1 U8505 ( .A(n12747), .B(n12780), .C(n4425), .Y(n8522) );
  NAND2X1 U8506 ( .A(ram[4085]), .B(n12780), .Y(n4425) );
  OAI21X1 U8507 ( .A(n12741), .B(n12780), .C(n4426), .Y(n8523) );
  NAND2X1 U8508 ( .A(ram[4086]), .B(n12780), .Y(n4426) );
  OAI21X1 U8509 ( .A(n12735), .B(n12780), .C(n4427), .Y(n8524) );
  NAND2X1 U8510 ( .A(ram[4087]), .B(n12780), .Y(n4427) );
  OAI21X1 U8511 ( .A(n12729), .B(n12780), .C(n4428), .Y(n8525) );
  NAND2X1 U8512 ( .A(ram[4088]), .B(n12780), .Y(n4428) );
  OAI21X1 U8513 ( .A(n12723), .B(n12780), .C(n4429), .Y(n8526) );
  NAND2X1 U8514 ( .A(ram[4089]), .B(n12780), .Y(n4429) );
  OAI21X1 U8515 ( .A(n12717), .B(n12780), .C(n4430), .Y(n8527) );
  NAND2X1 U8516 ( .A(ram[4090]), .B(n12780), .Y(n4430) );
  OAI21X1 U8517 ( .A(n12711), .B(n12780), .C(n4431), .Y(n8528) );
  NAND2X1 U8518 ( .A(ram[4091]), .B(n12780), .Y(n4431) );
  OAI21X1 U8519 ( .A(n12705), .B(n12780), .C(n4432), .Y(n8529) );
  NAND2X1 U8520 ( .A(ram[4092]), .B(n12780), .Y(n4432) );
  OAI21X1 U8521 ( .A(n12699), .B(n12780), .C(n4433), .Y(n8530) );
  NAND2X1 U8522 ( .A(ram[4093]), .B(n12780), .Y(n4433) );
  OAI21X1 U8523 ( .A(n12695), .B(n12780), .C(n4434), .Y(n8531) );
  NAND2X1 U8524 ( .A(ram[4094]), .B(n12780), .Y(n4434) );
  OAI21X1 U8525 ( .A(n12689), .B(n12780), .C(n4435), .Y(n8532) );
  NAND2X1 U8526 ( .A(ram[4095]), .B(n12780), .Y(n4435) );
  AND2X1 U8529 ( .A(mem_access_addr[1]), .B(mem_access_addr[0]), .Y(n4228) );
  AND2X1 U8530 ( .A(mem_access_addr[3]), .B(mem_access_addr[2]), .Y(n4384) );
  NAND3X1 U8531 ( .A(n1149), .B(mem_write_en), .C(n3609), .Y(n4436) );
  AND2X1 U8532 ( .A(mem_access_addr[7]), .B(mem_access_addr[6]), .Y(n3609) );
  AND2X1 U8533 ( .A(mem_access_addr[5]), .B(mem_access_addr[4]), .Y(n1149) );
  INVX1 U2 ( .A(n13039), .Y(n1) );
  INVX1 U3 ( .A(mem_access_addr[6]), .Y(n13039) );
  BUFX2 U4 ( .A(n12635), .Y(n12649) );
  BUFX2 U5 ( .A(n12635), .Y(n12648) );
  BUFX2 U6 ( .A(n12634), .Y(n12653) );
  BUFX2 U7 ( .A(n12634), .Y(n12654) );
  BUFX2 U8 ( .A(n12635), .Y(n12650) );
  BUFX2 U9 ( .A(n12634), .Y(n12652) );
  BUFX2 U10 ( .A(n12635), .Y(n12651) );
  BUFX2 U11 ( .A(n12632), .Y(n12658) );
  BUFX2 U12 ( .A(n12632), .Y(n12659) );
  BUFX2 U13 ( .A(n12633), .Y(n12655) );
  BUFX2 U14 ( .A(n12633), .Y(n12656) );
  BUFX2 U15 ( .A(n12633), .Y(n12657) );
  BUFX2 U16 ( .A(n12630), .Y(n12664) );
  BUFX2 U17 ( .A(n12630), .Y(n12665) );
  BUFX2 U18 ( .A(n12632), .Y(n12660) );
  BUFX2 U19 ( .A(n12631), .Y(n12661) );
  BUFX2 U20 ( .A(n12631), .Y(n12663) );
  BUFX2 U21 ( .A(n12631), .Y(n12662) );
  BUFX2 U22 ( .A(n12629), .Y(n12669) );
  BUFX2 U23 ( .A(n12628), .Y(n12670) );
  BUFX2 U24 ( .A(n12630), .Y(n12666) );
  BUFX2 U25 ( .A(n12629), .Y(n12667) );
  BUFX2 U26 ( .A(n12629), .Y(n12668) );
  BUFX2 U27 ( .A(n12627), .Y(n12674) );
  BUFX2 U28 ( .A(n12627), .Y(n12675) );
  BUFX2 U29 ( .A(n12628), .Y(n12671) );
  BUFX2 U30 ( .A(n12628), .Y(n12672) );
  BUFX2 U31 ( .A(n12627), .Y(n12673) );
  BUFX2 U32 ( .A(n12625), .Y(n12680) );
  BUFX2 U33 ( .A(n12625), .Y(n12681) );
  BUFX2 U34 ( .A(n12626), .Y(n12676) );
  BUFX2 U35 ( .A(n12626), .Y(n12677) );
  BUFX2 U36 ( .A(n12626), .Y(n12678) );
  BUFX2 U37 ( .A(n12625), .Y(n12679) );
  BUFX2 U70 ( .A(n12636), .Y(n12645) );
  BUFX2 U103 ( .A(n12636), .Y(n12646) );
  BUFX2 U136 ( .A(n12636), .Y(n12647) );
  BUFX2 U169 ( .A(n12637), .Y(n12642) );
  BUFX2 U202 ( .A(n12637), .Y(n12644) );
  BUFX2 U235 ( .A(n12637), .Y(n12643) );
  BUFX2 U268 ( .A(n12638), .Y(n12640) );
  BUFX2 U301 ( .A(n12638), .Y(n12641) );
  BUFX2 U334 ( .A(n12586), .Y(n12575) );
  BUFX2 U367 ( .A(n12588), .Y(n12576) );
  BUFX2 U400 ( .A(n12587), .Y(n12577) );
  BUFX2 U433 ( .A(n12587), .Y(n12578) );
  BUFX2 U466 ( .A(n12587), .Y(n12579) );
  BUFX2 U499 ( .A(n12588), .Y(n12580) );
  BUFX2 U532 ( .A(n12588), .Y(n12581) );
  BUFX2 U565 ( .A(n12588), .Y(n12582) );
  BUFX2 U599 ( .A(n12589), .Y(n12583) );
  BUFX2 U632 ( .A(n12589), .Y(n12584) );
  BUFX2 U665 ( .A(n12589), .Y(n12585) );
  BUFX2 U698 ( .A(n12638), .Y(n12639) );
  BUFX2 U731 ( .A(mem_access_addr[0]), .Y(n12634) );
  BUFX2 U764 ( .A(n12683), .Y(n12635) );
  BUFX2 U797 ( .A(n12622), .Y(n12633) );
  BUFX2 U830 ( .A(n12622), .Y(n12632) );
  BUFX2 U863 ( .A(n12622), .Y(n12631) );
  BUFX2 U896 ( .A(n12623), .Y(n12630) );
  BUFX2 U929 ( .A(n12623), .Y(n12629) );
  BUFX2 U962 ( .A(n12623), .Y(n12628) );
  BUFX2 U995 ( .A(n12624), .Y(n12627) );
  BUFX2 U1028 ( .A(n12624), .Y(n12626) );
  BUFX2 U1061 ( .A(n12624), .Y(n12625) );
  BUFX2 U1094 ( .A(n12595), .Y(n12597) );
  BUFX2 U1128 ( .A(n12596), .Y(n12598) );
  BUFX2 U1161 ( .A(n12595), .Y(n12601) );
  BUFX2 U1194 ( .A(n12596), .Y(n12599) );
  BUFX2 U1227 ( .A(n12596), .Y(n12600) );
  BUFX2 U1260 ( .A(n12595), .Y(n12603) );
  BUFX2 U1293 ( .A(n12595), .Y(n12602) );
  BUFX2 U1326 ( .A(n12594), .Y(n12606) );
  BUFX2 U1359 ( .A(n12594), .Y(n12604) );
  BUFX2 U1392 ( .A(n12594), .Y(n12605) );
  BUFX2 U1425 ( .A(n12593), .Y(n12609) );
  BUFX2 U1458 ( .A(n12593), .Y(n12607) );
  BUFX2 U1491 ( .A(n12593), .Y(n12608) );
  BUFX2 U1524 ( .A(n12592), .Y(n12610) );
  BUFX2 U1557 ( .A(n12592), .Y(n12611) );
  BUFX2 U1590 ( .A(n12591), .Y(n12614) );
  BUFX2 U1623 ( .A(n12592), .Y(n12612) );
  BUFX2 U1657 ( .A(n12591), .Y(n12613) );
  BUFX2 U1690 ( .A(n12591), .Y(n12615) );
  BUFX2 U1723 ( .A(n12590), .Y(n12617) );
  BUFX2 U1756 ( .A(n12590), .Y(n12616) );
  BUFX2 U1789 ( .A(n12683), .Y(n12622) );
  BUFX2 U1822 ( .A(n12683), .Y(n12623) );
  BUFX2 U1855 ( .A(n12683), .Y(n12624) );
  BUFX2 U1888 ( .A(n12586), .Y(n12587) );
  BUFX2 U1921 ( .A(n12586), .Y(n12588) );
  BUFX2 U1954 ( .A(n12586), .Y(n12589) );
  BUFX2 U1987 ( .A(n12621), .Y(n12636) );
  BUFX2 U2020 ( .A(n12621), .Y(n12637) );
  BUFX2 U2053 ( .A(n12621), .Y(n12638) );
  INVX2 U2086 ( .A(n3627), .Y(n13034) );
  INVX2 U2119 ( .A(n3644), .Y(n13033) );
  INVX2 U2152 ( .A(n3661), .Y(n13032) );
  INVX2 U2187 ( .A(n3678), .Y(n13031) );
  INVX2 U2220 ( .A(n3695), .Y(n13030) );
  INVX2 U2253 ( .A(n2), .Y(n13029) );
  INVX2 U2286 ( .A(n3780), .Y(n13028) );
  INVX2 U2319 ( .A(n3712), .Y(n13027) );
  INVX2 U2352 ( .A(n3729), .Y(n13026) );
  INVX2 U2385 ( .A(n3), .Y(n13025) );
  INVX2 U2418 ( .A(n3797), .Y(n13024) );
  INVX2 U2451 ( .A(n3746), .Y(n13023) );
  INVX2 U2484 ( .A(n3763), .Y(n13022) );
  INVX2 U2517 ( .A(n4), .Y(n13021) );
  INVX2 U2550 ( .A(n3814), .Y(n13020) );
  INVX2 U2583 ( .A(n31), .Y(n13019) );
  INVX2 U2616 ( .A(n32), .Y(n13018) );
  INVX2 U2649 ( .A(n33), .Y(n13017) );
  INVX2 U2682 ( .A(n34), .Y(n13016) );
  INVX2 U2716 ( .A(n24), .Y(n13015) );
  INVX2 U2749 ( .A(n35), .Y(n13014) );
  INVX2 U2782 ( .A(n55), .Y(n13013) );
  INVX2 U2815 ( .A(n73), .Y(n13012) );
  INVX2 U2848 ( .A(n91), .Y(n13011) );
  INVX2 U2881 ( .A(n36), .Y(n13010) );
  INVX2 U2914 ( .A(n109), .Y(n13009) );
  INVX2 U2947 ( .A(n127), .Y(n13008) );
  INVX2 U2980 ( .A(n25), .Y(n13007) );
  INVX2 U3013 ( .A(n37), .Y(n13006) );
  INVX2 U3046 ( .A(n145), .Y(n13005) );
  INVX2 U3079 ( .A(n163), .Y(n13004) );
  INVX2 U3112 ( .A(n181), .Y(n13003) );
  INVX2 U3145 ( .A(n199), .Y(n13002) );
  INVX2 U3178 ( .A(n217), .Y(n13001) );
  INVX2 U3211 ( .A(n235), .Y(n13000) );
  INVX2 U3245 ( .A(n253), .Y(n12999) );
  INVX2 U3278 ( .A(n271), .Y(n12998) );
  INVX2 U3311 ( .A(n345), .Y(n12997) );
  INVX2 U3344 ( .A(n362), .Y(n12996) );
  INVX2 U3377 ( .A(n289), .Y(n12995) );
  INVX2 U3410 ( .A(n307), .Y(n12994) );
  INVX2 U3443 ( .A(n379), .Y(n12993) );
  INVX2 U3476 ( .A(n396), .Y(n12992) );
  INVX2 U3509 ( .A(n26), .Y(n12991) );
  INVX2 U3542 ( .A(n328), .Y(n12990) );
  INVX2 U3575 ( .A(n413), .Y(n12989) );
  INVX2 U3608 ( .A(n430), .Y(n12988) );
  INVX2 U3641 ( .A(n447), .Y(n12987) );
  INVX2 U3674 ( .A(n464), .Y(n12986) );
  INVX2 U3707 ( .A(n481), .Y(n12985) );
  INVX2 U3740 ( .A(n498), .Y(n12984) );
  INVX2 U3774 ( .A(n515), .Y(n12983) );
  INVX2 U3807 ( .A(n532), .Y(n12982) );
  INVX2 U3840 ( .A(n583), .Y(n12981) );
  INVX2 U3873 ( .A(n602), .Y(n12980) );
  INVX2 U3906 ( .A(n549), .Y(n12979) );
  INVX2 U3939 ( .A(n566), .Y(n12978) );
  INVX2 U3972 ( .A(n653), .Y(n12977) );
  INVX2 U4005 ( .A(n670), .Y(n12976) );
  INVX2 U4038 ( .A(n619), .Y(n12975) );
  INVX2 U4071 ( .A(n636), .Y(n12974) );
  INVX2 U4104 ( .A(n687), .Y(n12973) );
  INVX2 U4137 ( .A(n704), .Y(n12972) );
  INVX2 U4170 ( .A(n721), .Y(n12971) );
  INVX2 U4203 ( .A(n738), .Y(n12970) );
  INVX2 U4236 ( .A(n755), .Y(n12969) );
  INVX2 U4269 ( .A(n772), .Y(n12968) );
  INVX2 U4304 ( .A(n27), .Y(n12967) );
  INVX2 U4337 ( .A(n789), .Y(n12966) );
  INVX2 U4370 ( .A(n857), .Y(n12965) );
  INVX2 U4403 ( .A(n876), .Y(n12964) );
  INVX2 U4436 ( .A(n806), .Y(n12963) );
  INVX2 U4469 ( .A(n823), .Y(n12962) );
  INVX2 U4502 ( .A(n893), .Y(n12961) );
  INVX2 U4535 ( .A(n910), .Y(n12960) );
  INVX2 U4568 ( .A(n28), .Y(n12959) );
  INVX2 U4601 ( .A(n840), .Y(n12958) );
  INVX2 U4634 ( .A(n927), .Y(n12957) );
  INVX2 U4667 ( .A(n944), .Y(n12956) );
  INVX2 U4700 ( .A(n5), .Y(n12955) );
  INVX2 U4733 ( .A(n6), .Y(n12954) );
  INVX2 U4766 ( .A(n961), .Y(n12953) );
  INVX2 U4799 ( .A(n978), .Y(n12952) );
  INVX2 U4833 ( .A(n7), .Y(n12951) );
  INVX2 U4866 ( .A(n8), .Y(n12950) );
  INVX2 U4899 ( .A(n1012), .Y(n12949) );
  INVX2 U4932 ( .A(n9), .Y(n12948) );
  INVX2 U4965 ( .A(n1029), .Y(n12947) );
  INVX2 U4998 ( .A(n995), .Y(n12946) );
  INVX2 U5031 ( .A(n1046), .Y(n12945) );
  INVX2 U5064 ( .A(n10), .Y(n12944) );
  INVX2 U5097 ( .A(n11), .Y(n12943) );
  INVX2 U5130 ( .A(n12), .Y(n12942) );
  INVX2 U5163 ( .A(n1063), .Y(n12941) );
  INVX2 U5196 ( .A(n13), .Y(n12940) );
  INVX2 U5229 ( .A(n1080), .Y(n12939) );
  INVX2 U5262 ( .A(n1097), .Y(n12938) );
  INVX2 U5295 ( .A(n1114), .Y(n12937) );
  INVX2 U5328 ( .A(n1131), .Y(n12936) );
  INVX2 U5362 ( .A(n1150), .Y(n12935) );
  INVX2 U5395 ( .A(n1167), .Y(n12934) );
  INVX2 U5428 ( .A(n1201), .Y(n12933) );
  INVX2 U5461 ( .A(n1218), .Y(n12932) );
  INVX2 U5494 ( .A(n1235), .Y(n12931) );
  INVX2 U5527 ( .A(n1252), .Y(n12930) );
  INVX2 U5560 ( .A(n1269), .Y(n12929) );
  INVX2 U5593 ( .A(n1286), .Y(n12928) );
  INVX2 U5626 ( .A(n1303), .Y(n12927) );
  INVX2 U5659 ( .A(n1184), .Y(n12926) );
  INVX2 U5692 ( .A(n1320), .Y(n12925) );
  INVX2 U5725 ( .A(n1337), .Y(n12924) );
  INVX2 U5758 ( .A(n1354), .Y(n12923) );
  INVX2 U5791 ( .A(n1371), .Y(n12922) );
  INVX2 U5824 ( .A(n1388), .Y(n12921) );
  INVX2 U5857 ( .A(n1405), .Y(n12920) );
  INVX2 U5891 ( .A(n1424), .Y(n12919) );
  INVX2 U5924 ( .A(n1441), .Y(n12918) );
  INVX2 U5957 ( .A(n1475), .Y(n12917) );
  INVX2 U5990 ( .A(n1492), .Y(n12916) );
  INVX2 U6023 ( .A(n1509), .Y(n12915) );
  INVX2 U6056 ( .A(n1526), .Y(n12914) );
  INVX2 U6089 ( .A(n1543), .Y(n12913) );
  INVX2 U6122 ( .A(n1560), .Y(n12912) );
  INVX2 U6155 ( .A(n1577), .Y(n12911) );
  INVX2 U6188 ( .A(n1458), .Y(n12910) );
  INVX2 U6221 ( .A(n1594), .Y(n12909) );
  INVX2 U6254 ( .A(n1611), .Y(n12908) );
  INVX2 U6287 ( .A(n1628), .Y(n12907) );
  INVX2 U6320 ( .A(n1645), .Y(n12906) );
  INVX2 U6353 ( .A(n1662), .Y(n12905) );
  INVX2 U6386 ( .A(n1679), .Y(n12904) );
  INVX2 U6421 ( .A(n1697), .Y(n12903) );
  INVX2 U6454 ( .A(n1714), .Y(n12902) );
  INVX2 U6487 ( .A(n1782), .Y(n12901) );
  INVX2 U6520 ( .A(n1799), .Y(n12900) );
  INVX2 U6553 ( .A(n1731), .Y(n12899) );
  INVX2 U6586 ( .A(n1748), .Y(n12898) );
  INVX2 U6619 ( .A(n1816), .Y(n12897) );
  INVX2 U6652 ( .A(n1833), .Y(n12896) );
  INVX2 U6685 ( .A(n29), .Y(n12895) );
  INVX2 U6718 ( .A(n1765), .Y(n12894) );
  INVX2 U6751 ( .A(n1850), .Y(n12893) );
  INVX2 U6784 ( .A(n1867), .Y(n12892) );
  INVX2 U6817 ( .A(n1884), .Y(n12891) );
  INVX2 U6850 ( .A(n1901), .Y(n12890) );
  INVX2 U6883 ( .A(n1918), .Y(n12889) );
  INVX2 U6916 ( .A(n1935), .Y(n12888) );
  INVX2 U6951 ( .A(n1952), .Y(n12887) );
  INVX2 U6984 ( .A(n1970), .Y(n12886) );
  INVX2 U7017 ( .A(n2004), .Y(n12885) );
  INVX2 U7050 ( .A(n14), .Y(n12884) );
  INVX2 U7083 ( .A(n2021), .Y(n12883) );
  INVX2 U7116 ( .A(n1987), .Y(n12882) );
  INVX2 U7149 ( .A(n2038), .Y(n12881) );
  INVX2 U7182 ( .A(n15), .Y(n12880) );
  INVX2 U7215 ( .A(n16), .Y(n12879) );
  INVX2 U7248 ( .A(n17), .Y(n12878) );
  INVX2 U7281 ( .A(n2055), .Y(n12877) );
  INVX2 U7314 ( .A(n18), .Y(n12876) );
  INVX2 U7347 ( .A(n2072), .Y(n12875) );
  INVX2 U7380 ( .A(n2089), .Y(n12874) );
  INVX2 U7413 ( .A(n2106), .Y(n12873) );
  INVX2 U7446 ( .A(n2123), .Y(n12872) );
  INVX2 U7481 ( .A(n2140), .Y(n12871) );
  INVX2 U7514 ( .A(n2157), .Y(n12870) );
  INVX2 U7547 ( .A(n2191), .Y(n12869) );
  INVX2 U7580 ( .A(n2208), .Y(n12868) );
  INVX2 U7613 ( .A(n2225), .Y(n12867) );
  INVX2 U7646 ( .A(n2243), .Y(n12866) );
  INVX2 U7679 ( .A(n2260), .Y(n12865) );
  INVX2 U7712 ( .A(n2277), .Y(n12864) );
  INVX2 U7745 ( .A(n2294), .Y(n12863) );
  INVX2 U7778 ( .A(n2174), .Y(n12862) );
  INVX2 U7811 ( .A(n2311), .Y(n12861) );
  INVX2 U7844 ( .A(n2328), .Y(n12860) );
  INVX2 U7877 ( .A(n2345), .Y(n12859) );
  INVX2 U7910 ( .A(n2362), .Y(n12858) );
  INVX2 U7943 ( .A(n2379), .Y(n12857) );
  INVX2 U7976 ( .A(n2396), .Y(n12856) );
  INVX2 U8011 ( .A(n2413), .Y(n12855) );
  INVX2 U8012 ( .A(n2430), .Y(n12854) );
  INVX2 U8045 ( .A(n2464), .Y(n12853) );
  INVX2 U8046 ( .A(n2481), .Y(n12852) );
  INVX2 U8079 ( .A(n2498), .Y(n12851) );
  INVX2 U8080 ( .A(n2517), .Y(n12850) );
  INVX2 U8113 ( .A(n2534), .Y(n12849) );
  INVX2 U8114 ( .A(n2551), .Y(n12848) );
  INVX2 U8148 ( .A(n2568), .Y(n12847) );
  INVX2 U8149 ( .A(n2447), .Y(n12846) );
  INVX2 U8182 ( .A(n2585), .Y(n12845) );
  INVX2 U8183 ( .A(n2602), .Y(n12844) );
  INVX2 U8216 ( .A(n2619), .Y(n12843) );
  INVX2 U8217 ( .A(n2636), .Y(n12842) );
  INVX2 U8250 ( .A(n2653), .Y(n12841) );
  INVX2 U8251 ( .A(n2670), .Y(n12840) );
  INVX2 U8285 ( .A(n2687), .Y(n12839) );
  INVX2 U8286 ( .A(n2704), .Y(n12838) );
  INVX2 U8319 ( .A(n2772), .Y(n12837) );
  INVX2 U8320 ( .A(n2790), .Y(n12836) );
  INVX2 U8353 ( .A(n2721), .Y(n12835) );
  INVX2 U8354 ( .A(n2738), .Y(n12834) );
  INVX2 U8387 ( .A(n2807), .Y(n12833) );
  INVX2 U8388 ( .A(n2824), .Y(n12832) );
  INVX2 U8422 ( .A(n30), .Y(n12831) );
  INVX2 U8423 ( .A(n2755), .Y(n12830) );
  INVX2 U8457 ( .A(n2841), .Y(n12829) );
  INVX2 U8458 ( .A(n2858), .Y(n12828) );
  INVX2 U8492 ( .A(n2875), .Y(n12827) );
  INVX2 U8493 ( .A(n2892), .Y(n12826) );
  INVX2 U8527 ( .A(n2909), .Y(n12825) );
  INVX2 U8528 ( .A(n2926), .Y(n12824) );
  INVX2 U8534 ( .A(n2943), .Y(n12823) );
  INVX2 U8535 ( .A(n2960), .Y(n12822) );
  INVX2 U8536 ( .A(n2994), .Y(n12821) );
  INVX2 U8537 ( .A(n19), .Y(n12820) );
  INVX2 U8538 ( .A(n3011), .Y(n12819) );
  INVX2 U8539 ( .A(n2977), .Y(n12818) );
  INVX2 U8540 ( .A(n3028), .Y(n12817) );
  INVX2 U8541 ( .A(n20), .Y(n12816) );
  INVX2 U8542 ( .A(n21), .Y(n12815) );
  INVX2 U8543 ( .A(n22), .Y(n12814) );
  INVX2 U8544 ( .A(n3045), .Y(n12813) );
  INVX2 U8545 ( .A(n23), .Y(n12812) );
  INVX2 U8546 ( .A(n3063), .Y(n12811) );
  INVX2 U8547 ( .A(n3080), .Y(n12810) );
  INVX2 U8548 ( .A(n3097), .Y(n12809) );
  INVX2 U8549 ( .A(n3114), .Y(n12808) );
  INVX2 U8550 ( .A(n3131), .Y(n12807) );
  INVX2 U8551 ( .A(n3148), .Y(n12806) );
  INVX2 U8552 ( .A(n3182), .Y(n12805) );
  INVX2 U8553 ( .A(n3199), .Y(n12804) );
  INVX2 U8554 ( .A(n3216), .Y(n12803) );
  INVX2 U8555 ( .A(n3233), .Y(n12802) );
  INVX2 U8556 ( .A(n3250), .Y(n12801) );
  INVX2 U8557 ( .A(n3267), .Y(n12800) );
  INVX2 U8558 ( .A(n3284), .Y(n12799) );
  INVX2 U8559 ( .A(n3165), .Y(n12798) );
  INVX2 U8560 ( .A(n3301), .Y(n12797) );
  INVX2 U8561 ( .A(n3318), .Y(n12796) );
  INVX2 U8562 ( .A(n3336), .Y(n12795) );
  INVX2 U8563 ( .A(n3353), .Y(n12794) );
  INVX2 U8564 ( .A(n3370), .Y(n12793) );
  INVX2 U8565 ( .A(n3387), .Y(n12792) );
  INVX2 U8566 ( .A(n3404), .Y(n12791) );
  INVX2 U8567 ( .A(n3421), .Y(n12790) );
  INVX2 U8568 ( .A(n3472), .Y(n12789) );
  INVX2 U8569 ( .A(n3489), .Y(n12788) );
  INVX2 U8570 ( .A(n3506), .Y(n12787) );
  INVX2 U8571 ( .A(n3438), .Y(n12786) );
  INVX2 U8572 ( .A(n3523), .Y(n12785) );
  INVX2 U8573 ( .A(n3540), .Y(n12784) );
  INVX2 U8574 ( .A(n3557), .Y(n12783) );
  INVX2 U8575 ( .A(n3455), .Y(n12782) );
  INVX2 U8576 ( .A(n3574), .Y(n12781) );
  INVX2 U8577 ( .A(n3591), .Y(n12780) );
  INVX2 U8578 ( .A(n3610), .Y(n13035) );
  BUFX2 U8579 ( .A(n12620), .Y(n12596) );
  BUFX2 U8580 ( .A(n12620), .Y(n12595) );
  BUFX2 U8581 ( .A(n12619), .Y(n12594) );
  BUFX2 U8582 ( .A(n12619), .Y(n12593) );
  BUFX2 U8583 ( .A(n12619), .Y(n12592) );
  BUFX2 U8584 ( .A(mem_access_addr[0]), .Y(n12683) );
  BUFX2 U8585 ( .A(n12618), .Y(n12591) );
  BUFX2 U8586 ( .A(mem_access_addr[2]), .Y(n12586) );
  BUFX2 U8587 ( .A(n12682), .Y(n12621) );
  BUFX2 U8588 ( .A(mem_access_addr[0]), .Y(n12682) );
  BUFX2 U8589 ( .A(n12618), .Y(n12590) );
  AND2X1 U8590 ( .A(n162), .B(n13043), .Y(n2) );
  AND2X1 U8591 ( .A(n234), .B(n13043), .Y(n3) );
  AND2X1 U8592 ( .A(n306), .B(n13043), .Y(n4) );
  AND2X1 U8593 ( .A(n13046), .B(n54), .Y(n5) );
  AND2X1 U8594 ( .A(n13046), .B(n72), .Y(n6) );
  AND2X1 U8595 ( .A(n13046), .B(n126), .Y(n7) );
  AND2X1 U8596 ( .A(n13046), .B(n144), .Y(n8) );
  AND2X1 U8597 ( .A(n13046), .B(n180), .Y(n9) );
  AND2X1 U8598 ( .A(n13046), .B(n252), .Y(n10) );
  AND2X1 U8599 ( .A(n13046), .B(n270), .Y(n11) );
  AND2X1 U8600 ( .A(n13046), .B(n288), .Y(n12) );
  AND2X1 U8601 ( .A(n13046), .B(n324), .Y(n13) );
  AND2X1 U8602 ( .A(n13050), .B(n180), .Y(n14) );
  AND2X1 U8603 ( .A(n13050), .B(n252), .Y(n15) );
  AND2X1 U8604 ( .A(n13050), .B(n270), .Y(n16) );
  AND2X1 U8605 ( .A(n13050), .B(n288), .Y(n17) );
  AND2X1 U8606 ( .A(n13050), .B(n324), .Y(n18) );
  AND2X1 U8607 ( .A(n13054), .B(n180), .Y(n19) );
  AND2X1 U8608 ( .A(n13054), .B(n252), .Y(n20) );
  AND2X1 U8609 ( .A(n13054), .B(n270), .Y(n21) );
  AND2X1 U8610 ( .A(n13054), .B(n288), .Y(n22) );
  AND2X1 U8611 ( .A(n13054), .B(n324), .Y(n23) );
  AND2X1 U8612 ( .A(n13042), .B(n126), .Y(n24) );
  AND2X1 U8613 ( .A(n13042), .B(n270), .Y(n25) );
  AND2X1 U8614 ( .A(n13041), .B(n270), .Y(n26) );
  AND2X1 U8615 ( .A(n13047), .B(n126), .Y(n27) );
  AND2X1 U8616 ( .A(n13047), .B(n270), .Y(n28) );
  AND2X1 U8617 ( .A(n13051), .B(n270), .Y(n29) );
  AND2X1 U8618 ( .A(n13055), .B(n270), .Y(n30) );
  BUFX2 U8619 ( .A(mem_access_addr[4]), .Y(n12565) );
  BUFX2 U8620 ( .A(mem_access_addr[4]), .Y(n12566) );
  BUFX2 U8621 ( .A(mem_access_addr[4]), .Y(n12567) );
  BUFX2 U8622 ( .A(mem_access_addr[3]), .Y(n12568) );
  BUFX2 U8623 ( .A(n12574), .Y(n12569) );
  BUFX2 U8624 ( .A(n12574), .Y(n12570) );
  BUFX2 U8625 ( .A(n12574), .Y(n12571) );
  BUFX2 U8626 ( .A(n12574), .Y(n12572) );
  BUFX2 U8627 ( .A(mem_access_addr[3]), .Y(n12573) );
  BUFX2 U8628 ( .A(n12775), .Y(n12776) );
  BUFX2 U8629 ( .A(n12769), .Y(n12770) );
  BUFX2 U8630 ( .A(n12763), .Y(n12764) );
  BUFX2 U8631 ( .A(n12757), .Y(n12758) );
  BUFX2 U8632 ( .A(n12751), .Y(n12752) );
  BUFX2 U8633 ( .A(n12745), .Y(n12746) );
  BUFX2 U8634 ( .A(n12739), .Y(n12740) );
  BUFX2 U8635 ( .A(n12733), .Y(n12734) );
  BUFX2 U8636 ( .A(n12727), .Y(n12728) );
  BUFX2 U8637 ( .A(n12721), .Y(n12722) );
  BUFX2 U8638 ( .A(n12715), .Y(n12716) );
  BUFX2 U8639 ( .A(n12709), .Y(n12710) );
  BUFX2 U8640 ( .A(n12703), .Y(n12704) );
  BUFX2 U8641 ( .A(n12697), .Y(n12698) );
  BUFX2 U8642 ( .A(n12691), .Y(n12692) );
  BUFX2 U8643 ( .A(n12685), .Y(n12686) );
  BUFX2 U8644 ( .A(n12774), .Y(n12777) );
  BUFX2 U8645 ( .A(n12768), .Y(n12771) );
  BUFX2 U8646 ( .A(n12762), .Y(n12765) );
  BUFX2 U8647 ( .A(n12756), .Y(n12759) );
  BUFX2 U8648 ( .A(n12750), .Y(n12753) );
  BUFX2 U8649 ( .A(n12744), .Y(n12747) );
  BUFX2 U8650 ( .A(n12738), .Y(n12741) );
  BUFX2 U8651 ( .A(n12732), .Y(n12735) );
  BUFX2 U8652 ( .A(n12726), .Y(n12729) );
  BUFX2 U8653 ( .A(n12720), .Y(n12723) );
  BUFX2 U8654 ( .A(n12714), .Y(n12717) );
  BUFX2 U8655 ( .A(n12708), .Y(n12711) );
  BUFX2 U8656 ( .A(n12702), .Y(n12705) );
  BUFX2 U8657 ( .A(n12696), .Y(n12699) );
  BUFX2 U8658 ( .A(n12690), .Y(n12693) );
  BUFX2 U8659 ( .A(n12684), .Y(n12687) );
  BUFX2 U8660 ( .A(n12774), .Y(n12778) );
  BUFX2 U8661 ( .A(n12768), .Y(n12772) );
  BUFX2 U8662 ( .A(n12762), .Y(n12766) );
  BUFX2 U8663 ( .A(n12756), .Y(n12760) );
  BUFX2 U8664 ( .A(n12750), .Y(n12754) );
  BUFX2 U8665 ( .A(n12744), .Y(n12748) );
  BUFX2 U8666 ( .A(n12738), .Y(n12742) );
  BUFX2 U8667 ( .A(n12732), .Y(n12736) );
  BUFX2 U8668 ( .A(n12726), .Y(n12730) );
  BUFX2 U8669 ( .A(n12720), .Y(n12724) );
  BUFX2 U8670 ( .A(n12714), .Y(n12718) );
  BUFX2 U8671 ( .A(n12708), .Y(n12712) );
  BUFX2 U8672 ( .A(n12702), .Y(n12706) );
  BUFX2 U8673 ( .A(n12696), .Y(n12700) );
  BUFX2 U8674 ( .A(n12690), .Y(n12694) );
  BUFX2 U8675 ( .A(n12684), .Y(n12688) );
  BUFX2 U8676 ( .A(n12774), .Y(n12779) );
  BUFX2 U8677 ( .A(n12768), .Y(n12773) );
  BUFX2 U8678 ( .A(n12762), .Y(n12767) );
  BUFX2 U8679 ( .A(n12756), .Y(n12761) );
  BUFX2 U8680 ( .A(n12750), .Y(n12755) );
  BUFX2 U8681 ( .A(n12744), .Y(n12749) );
  BUFX2 U8682 ( .A(n12738), .Y(n12743) );
  BUFX2 U8683 ( .A(n12732), .Y(n12737) );
  BUFX2 U8684 ( .A(n12726), .Y(n12731) );
  BUFX2 U8685 ( .A(n12720), .Y(n12725) );
  BUFX2 U8686 ( .A(n12714), .Y(n12719) );
  BUFX2 U8687 ( .A(n12708), .Y(n12713) );
  BUFX2 U8688 ( .A(n12702), .Y(n12707) );
  BUFX2 U8689 ( .A(n12696), .Y(n12701) );
  BUFX2 U8690 ( .A(n12690), .Y(n12695) );
  BUFX2 U8691 ( .A(n12684), .Y(n12689) );
  BUFX2 U8692 ( .A(mem_access_addr[4]), .Y(n12564) );
  AND2X1 U8693 ( .A(n13042), .B(n54), .Y(n31) );
  AND2X1 U8694 ( .A(n13042), .B(n72), .Y(n32) );
  AND2X1 U8695 ( .A(n13042), .B(n90), .Y(n33) );
  AND2X1 U8696 ( .A(n13042), .B(n108), .Y(n34) );
  AND2X1 U8697 ( .A(n13042), .B(n144), .Y(n35) );
  AND2X1 U8698 ( .A(n13042), .B(n216), .Y(n36) );
  AND2X1 U8699 ( .A(n13042), .B(n288), .Y(n37) );
  AND2X1 U8700 ( .A(n13042), .B(n162), .Y(n55) );
  AND2X1 U8701 ( .A(n13042), .B(n180), .Y(n73) );
  AND2X1 U8702 ( .A(n13042), .B(n198), .Y(n91) );
  AND2X1 U8703 ( .A(n13042), .B(n234), .Y(n109) );
  AND2X1 U8704 ( .A(n13042), .B(n252), .Y(n127) );
  AND2X1 U8705 ( .A(n13042), .B(n306), .Y(n145) );
  AND2X1 U8706 ( .A(n13042), .B(n324), .Y(n163) );
  AND2X1 U8707 ( .A(n13041), .B(n54), .Y(n181) );
  AND2X1 U8708 ( .A(n13041), .B(n72), .Y(n199) );
  AND2X1 U8709 ( .A(n13041), .B(n90), .Y(n217) );
  AND2X1 U8710 ( .A(n13041), .B(n108), .Y(n235) );
  AND2X1 U8711 ( .A(n13041), .B(n126), .Y(n253) );
  AND2X1 U8712 ( .A(n13041), .B(n144), .Y(n271) );
  AND2X1 U8713 ( .A(n13041), .B(n198), .Y(n289) );
  AND2X1 U8714 ( .A(n13041), .B(n216), .Y(n307) );
  AND2X1 U8715 ( .A(n13041), .B(n288), .Y(n328) );
  AND2X1 U8716 ( .A(n13041), .B(n162), .Y(n345) );
  AND2X1 U8717 ( .A(n13041), .B(n180), .Y(n362) );
  AND2X1 U8718 ( .A(n13041), .B(n234), .Y(n379) );
  AND2X1 U8719 ( .A(n13041), .B(n252), .Y(n396) );
  AND2X1 U8720 ( .A(n13041), .B(n306), .Y(n413) );
  AND2X1 U8721 ( .A(n13041), .B(n324), .Y(n430) );
  AND2X1 U8722 ( .A(n13040), .B(n54), .Y(n447) );
  AND2X1 U8723 ( .A(n13040), .B(n72), .Y(n464) );
  AND2X1 U8724 ( .A(n13040), .B(n90), .Y(n481) );
  AND2X1 U8725 ( .A(n13040), .B(n108), .Y(n498) );
  AND2X1 U8726 ( .A(n13040), .B(n126), .Y(n515) );
  AND2X1 U8727 ( .A(n13040), .B(n144), .Y(n532) );
  AND2X1 U8728 ( .A(n13040), .B(n198), .Y(n549) );
  AND2X1 U8729 ( .A(n13040), .B(n216), .Y(n566) );
  AND2X1 U8730 ( .A(n13040), .B(n162), .Y(n583) );
  AND2X1 U8731 ( .A(n13040), .B(n180), .Y(n602) );
  AND2X1 U8732 ( .A(n13040), .B(n270), .Y(n619) );
  AND2X1 U8733 ( .A(n13040), .B(n288), .Y(n636) );
  AND2X1 U8734 ( .A(n13040), .B(n234), .Y(n653) );
  AND2X1 U8735 ( .A(n13040), .B(n252), .Y(n670) );
  AND2X1 U8736 ( .A(n13040), .B(n306), .Y(n687) );
  AND2X1 U8737 ( .A(n13040), .B(n324), .Y(n704) );
  AND2X1 U8738 ( .A(n13047), .B(n54), .Y(n721) );
  AND2X1 U8739 ( .A(n13047), .B(n72), .Y(n738) );
  AND2X1 U8740 ( .A(n13047), .B(n90), .Y(n755) );
  AND2X1 U8741 ( .A(n13047), .B(n108), .Y(n772) );
  AND2X1 U8742 ( .A(n13047), .B(n144), .Y(n789) );
  AND2X1 U8743 ( .A(n13047), .B(n198), .Y(n806) );
  AND2X1 U8744 ( .A(n13047), .B(n216), .Y(n823) );
  AND2X1 U8745 ( .A(n13047), .B(n288), .Y(n840) );
  AND2X1 U8746 ( .A(n13047), .B(n162), .Y(n857) );
  AND2X1 U8747 ( .A(n13047), .B(n180), .Y(n876) );
  AND2X1 U8748 ( .A(n13047), .B(n234), .Y(n893) );
  AND2X1 U8749 ( .A(n13047), .B(n252), .Y(n910) );
  AND2X1 U8750 ( .A(n13047), .B(n306), .Y(n927) );
  AND2X1 U8751 ( .A(n13047), .B(n324), .Y(n944) );
  AND2X1 U8752 ( .A(n13046), .B(n90), .Y(n961) );
  AND2X1 U8753 ( .A(n13046), .B(n108), .Y(n978) );
  AND2X1 U8754 ( .A(n13046), .B(n216), .Y(n995) );
  AND2X1 U8755 ( .A(n13046), .B(n162), .Y(n1012) );
  AND2X1 U8756 ( .A(n13046), .B(n198), .Y(n1029) );
  AND2X1 U8757 ( .A(n13046), .B(n234), .Y(n1046) );
  AND2X1 U8758 ( .A(n13046), .B(n306), .Y(n1063) );
  AND2X1 U8759 ( .A(n13045), .B(n54), .Y(n1080) );
  AND2X1 U8760 ( .A(n13045), .B(n72), .Y(n1097) );
  AND2X1 U8761 ( .A(n13045), .B(n90), .Y(n1114) );
  AND2X1 U8762 ( .A(n13045), .B(n108), .Y(n1131) );
  AND2X1 U8763 ( .A(n13045), .B(n126), .Y(n1150) );
  AND2X1 U8764 ( .A(n13045), .B(n144), .Y(n1167) );
  AND2X1 U8765 ( .A(n13045), .B(n288), .Y(n1184) );
  AND2X1 U8766 ( .A(n13045), .B(n162), .Y(n1201) );
  AND2X1 U8767 ( .A(n13045), .B(n180), .Y(n1218) );
  AND2X1 U8768 ( .A(n13045), .B(n198), .Y(n1235) );
  AND2X1 U8769 ( .A(n13045), .B(n216), .Y(n1252) );
  AND2X1 U8770 ( .A(n13045), .B(n234), .Y(n1269) );
  AND2X1 U8771 ( .A(n13045), .B(n252), .Y(n1286) );
  AND2X1 U8772 ( .A(n13045), .B(n270), .Y(n1303) );
  AND2X1 U8773 ( .A(n13045), .B(n306), .Y(n1320) );
  AND2X1 U8774 ( .A(n13045), .B(n324), .Y(n1337) );
  AND2X1 U8775 ( .A(n13044), .B(n54), .Y(n1354) );
  AND2X1 U8776 ( .A(n13044), .B(n72), .Y(n1371) );
  AND2X1 U8777 ( .A(n13044), .B(n90), .Y(n1388) );
  AND2X1 U8778 ( .A(n13044), .B(n108), .Y(n1405) );
  AND2X1 U8779 ( .A(n13044), .B(n126), .Y(n1424) );
  AND2X1 U8780 ( .A(n13044), .B(n144), .Y(n1441) );
  AND2X1 U8781 ( .A(n13044), .B(n288), .Y(n1458) );
  AND2X1 U8782 ( .A(n13044), .B(n162), .Y(n1475) );
  AND2X1 U8783 ( .A(n13044), .B(n180), .Y(n1492) );
  AND2X1 U8784 ( .A(n13044), .B(n198), .Y(n1509) );
  AND2X1 U8785 ( .A(n13044), .B(n216), .Y(n1526) );
  AND2X1 U8786 ( .A(n13044), .B(n234), .Y(n1543) );
  AND2X1 U8787 ( .A(n13044), .B(n252), .Y(n1560) );
  AND2X1 U8788 ( .A(n13044), .B(n270), .Y(n1577) );
  AND2X1 U8789 ( .A(n13044), .B(n306), .Y(n1594) );
  AND2X1 U8790 ( .A(n13044), .B(n324), .Y(n1611) );
  AND2X1 U8791 ( .A(n13051), .B(n54), .Y(n1628) );
  AND2X1 U8792 ( .A(n13051), .B(n72), .Y(n1645) );
  AND2X1 U8793 ( .A(n13051), .B(n90), .Y(n1662) );
  AND2X1 U8794 ( .A(n13051), .B(n108), .Y(n1679) );
  AND2X1 U8795 ( .A(n13051), .B(n126), .Y(n1697) );
  AND2X1 U8796 ( .A(n13051), .B(n144), .Y(n1714) );
  AND2X1 U8797 ( .A(n13051), .B(n198), .Y(n1731) );
  AND2X1 U8798 ( .A(n13051), .B(n216), .Y(n1748) );
  AND2X1 U8799 ( .A(n13051), .B(n288), .Y(n1765) );
  AND2X1 U8800 ( .A(n13051), .B(n162), .Y(n1782) );
  AND2X1 U8801 ( .A(n13051), .B(n180), .Y(n1799) );
  AND2X1 U8802 ( .A(n13051), .B(n234), .Y(n1816) );
  AND2X1 U8803 ( .A(n13051), .B(n252), .Y(n1833) );
  AND2X1 U8804 ( .A(n13051), .B(n306), .Y(n1850) );
  AND2X1 U8805 ( .A(n13051), .B(n324), .Y(n1867) );
  AND2X1 U8806 ( .A(n13050), .B(n54), .Y(n1884) );
  AND2X1 U8807 ( .A(n13050), .B(n72), .Y(n1901) );
  AND2X1 U8808 ( .A(n13050), .B(n90), .Y(n1918) );
  AND2X1 U8809 ( .A(n13050), .B(n108), .Y(n1935) );
  AND2X1 U8810 ( .A(n13050), .B(n126), .Y(n1952) );
  AND2X1 U8811 ( .A(n13050), .B(n144), .Y(n1970) );
  AND2X1 U8812 ( .A(n13050), .B(n216), .Y(n1987) );
  AND2X1 U8813 ( .A(n13050), .B(n162), .Y(n2004) );
  AND2X1 U8814 ( .A(n13050), .B(n198), .Y(n2021) );
  AND2X1 U8815 ( .A(n13050), .B(n234), .Y(n2038) );
  AND2X1 U8816 ( .A(n13050), .B(n306), .Y(n2055) );
  AND2X1 U8817 ( .A(n13049), .B(n54), .Y(n2072) );
  AND2X1 U8818 ( .A(n13049), .B(n72), .Y(n2089) );
  AND2X1 U8819 ( .A(n13049), .B(n90), .Y(n2106) );
  AND2X1 U8820 ( .A(n13049), .B(n108), .Y(n2123) );
  AND2X1 U8821 ( .A(n13049), .B(n126), .Y(n2140) );
  AND2X1 U8822 ( .A(n13049), .B(n144), .Y(n2157) );
  AND2X1 U8823 ( .A(n13049), .B(n288), .Y(n2174) );
  AND2X1 U8824 ( .A(n13049), .B(n162), .Y(n2191) );
  AND2X1 U8825 ( .A(n13049), .B(n180), .Y(n2208) );
  AND2X1 U8826 ( .A(n13049), .B(n198), .Y(n2225) );
  AND2X1 U8827 ( .A(n13049), .B(n216), .Y(n2243) );
  AND2X1 U8828 ( .A(n13049), .B(n234), .Y(n2260) );
  AND2X1 U8829 ( .A(n13049), .B(n252), .Y(n2277) );
  AND2X1 U8830 ( .A(n13049), .B(n270), .Y(n2294) );
  AND2X1 U8831 ( .A(n13049), .B(n306), .Y(n2311) );
  AND2X1 U8832 ( .A(n13049), .B(n324), .Y(n2328) );
  AND2X1 U8833 ( .A(n13048), .B(n54), .Y(n2345) );
  AND2X1 U8834 ( .A(n13048), .B(n72), .Y(n2362) );
  AND2X1 U8835 ( .A(n13048), .B(n90), .Y(n2379) );
  AND2X1 U8836 ( .A(n13048), .B(n108), .Y(n2396) );
  AND2X1 U8837 ( .A(n13048), .B(n126), .Y(n2413) );
  AND2X1 U8838 ( .A(n13048), .B(n144), .Y(n2430) );
  AND2X1 U8839 ( .A(n13048), .B(n288), .Y(n2447) );
  AND2X1 U8840 ( .A(n13048), .B(n162), .Y(n2464) );
  AND2X1 U8841 ( .A(n13048), .B(n180), .Y(n2481) );
  AND2X1 U8842 ( .A(n13048), .B(n198), .Y(n2498) );
  AND2X1 U8843 ( .A(n13048), .B(n216), .Y(n2517) );
  AND2X1 U8844 ( .A(n13048), .B(n234), .Y(n2534) );
  AND2X1 U8845 ( .A(n13048), .B(n252), .Y(n2551) );
  AND2X1 U8846 ( .A(n13048), .B(n270), .Y(n2568) );
  AND2X1 U8847 ( .A(n13048), .B(n306), .Y(n2585) );
  AND2X1 U8848 ( .A(n13048), .B(n324), .Y(n2602) );
  AND2X1 U8849 ( .A(n13055), .B(n54), .Y(n2619) );
  AND2X1 U8850 ( .A(n13055), .B(n72), .Y(n2636) );
  AND2X1 U8851 ( .A(n13055), .B(n90), .Y(n2653) );
  AND2X1 U8852 ( .A(n13055), .B(n108), .Y(n2670) );
  AND2X1 U8853 ( .A(n13055), .B(n126), .Y(n2687) );
  AND2X1 U8854 ( .A(n13055), .B(n144), .Y(n2704) );
  AND2X1 U8855 ( .A(n13055), .B(n198), .Y(n2721) );
  AND2X1 U8856 ( .A(n13055), .B(n216), .Y(n2738) );
  AND2X1 U8857 ( .A(n13055), .B(n288), .Y(n2755) );
  AND2X1 U8858 ( .A(n13055), .B(n162), .Y(n2772) );
  AND2X1 U8859 ( .A(n13055), .B(n180), .Y(n2790) );
  AND2X1 U8860 ( .A(n13055), .B(n234), .Y(n2807) );
  AND2X1 U8861 ( .A(n13055), .B(n252), .Y(n2824) );
  AND2X1 U8862 ( .A(n13055), .B(n306), .Y(n2841) );
  AND2X1 U8863 ( .A(n13055), .B(n324), .Y(n2858) );
  AND2X1 U8864 ( .A(n13054), .B(n54), .Y(n2875) );
  AND2X1 U8865 ( .A(n13054), .B(n72), .Y(n2892) );
  AND2X1 U8866 ( .A(n13054), .B(n90), .Y(n2909) );
  AND2X1 U8867 ( .A(n13054), .B(n108), .Y(n2926) );
  AND2X1 U8868 ( .A(n13054), .B(n126), .Y(n2943) );
  AND2X1 U8869 ( .A(n13054), .B(n144), .Y(n2960) );
  AND2X1 U8870 ( .A(n13054), .B(n216), .Y(n2977) );
  AND2X1 U8871 ( .A(n13054), .B(n162), .Y(n2994) );
  AND2X1 U8872 ( .A(n13054), .B(n198), .Y(n3011) );
  AND2X1 U8873 ( .A(n13054), .B(n234), .Y(n3028) );
  AND2X1 U8874 ( .A(n13054), .B(n306), .Y(n3045) );
  AND2X1 U8875 ( .A(n13053), .B(n54), .Y(n3063) );
  AND2X1 U8876 ( .A(n13053), .B(n72), .Y(n3080) );
  AND2X1 U8877 ( .A(n13053), .B(n90), .Y(n3097) );
  AND2X1 U8878 ( .A(n13053), .B(n108), .Y(n3114) );
  AND2X1 U8879 ( .A(n13053), .B(n126), .Y(n3131) );
  AND2X1 U8880 ( .A(n13053), .B(n144), .Y(n3148) );
  AND2X1 U8881 ( .A(n13053), .B(n288), .Y(n3165) );
  AND2X1 U8882 ( .A(n13053), .B(n162), .Y(n3182) );
  AND2X1 U8883 ( .A(n13053), .B(n180), .Y(n3199) );
  AND2X1 U8884 ( .A(n13053), .B(n198), .Y(n3216) );
  AND2X1 U8885 ( .A(n13053), .B(n216), .Y(n3233) );
  AND2X1 U8886 ( .A(n13053), .B(n234), .Y(n3250) );
  AND2X1 U8887 ( .A(n13053), .B(n252), .Y(n3267) );
  AND2X1 U8888 ( .A(n13053), .B(n270), .Y(n3284) );
  AND2X1 U8889 ( .A(n13053), .B(n306), .Y(n3301) );
  AND2X1 U8890 ( .A(n13053), .B(n324), .Y(n3318) );
  AND2X1 U8891 ( .A(n13052), .B(n54), .Y(n3336) );
  AND2X1 U8892 ( .A(n13052), .B(n72), .Y(n3353) );
  AND2X1 U8893 ( .A(n13052), .B(n90), .Y(n3370) );
  AND2X1 U8894 ( .A(n13052), .B(n108), .Y(n3387) );
  AND2X1 U8895 ( .A(n13052), .B(n126), .Y(n3404) );
  AND2X1 U8896 ( .A(n13052), .B(n144), .Y(n3421) );
  AND2X1 U8897 ( .A(n13052), .B(n216), .Y(n3438) );
  AND2X1 U8898 ( .A(n13052), .B(n288), .Y(n3455) );
  AND2X1 U8899 ( .A(n13052), .B(n162), .Y(n3472) );
  AND2X1 U8900 ( .A(n13052), .B(n180), .Y(n3489) );
  AND2X1 U8901 ( .A(n13052), .B(n198), .Y(n3506) );
  AND2X1 U8902 ( .A(n13052), .B(n234), .Y(n3523) );
  AND2X1 U8903 ( .A(n13052), .B(n252), .Y(n3540) );
  AND2X1 U8904 ( .A(n13052), .B(n270), .Y(n3557) );
  AND2X1 U8905 ( .A(n13052), .B(n306), .Y(n3574) );
  AND2X1 U8906 ( .A(n13052), .B(n324), .Y(n3591) );
  AND2X1 U8907 ( .A(n54), .B(n13043), .Y(n3610) );
  AND2X1 U8908 ( .A(n72), .B(n13043), .Y(n3627) );
  AND2X1 U8909 ( .A(n90), .B(n13043), .Y(n3644) );
  AND2X1 U8910 ( .A(n108), .B(n13043), .Y(n3661) );
  AND2X1 U8911 ( .A(n126), .B(n13043), .Y(n3678) );
  AND2X1 U8912 ( .A(n144), .B(n13043), .Y(n3695) );
  AND2X1 U8913 ( .A(n198), .B(n13043), .Y(n3712) );
  AND2X1 U8914 ( .A(n216), .B(n13043), .Y(n3729) );
  AND2X1 U8915 ( .A(n270), .B(n13043), .Y(n3746) );
  AND2X1 U8916 ( .A(n288), .B(n13043), .Y(n3763) );
  AND2X1 U8917 ( .A(n180), .B(n13043), .Y(n3780) );
  AND2X1 U8918 ( .A(n252), .B(n13043), .Y(n3797) );
  AND2X1 U8919 ( .A(n324), .B(n13043), .Y(n3814) );
  BUFX2 U8920 ( .A(mem_access_addr[1]), .Y(n12620) );
  BUFX2 U8921 ( .A(mem_access_addr[1]), .Y(n12619) );
  BUFX2 U8922 ( .A(mem_access_addr[1]), .Y(n12618) );
  INVX2 U8923 ( .A(n2789), .Y(n13050) );
  INVX2 U8924 ( .A(n1148), .Y(n13040) );
  INVX2 U8925 ( .A(n1422), .Y(n13047) );
  INVX2 U8926 ( .A(n325), .Y(n13043) );
  INVX2 U8927 ( .A(n1696), .Y(n13046) );
  INVX2 U8928 ( .A(n1969), .Y(n13045) );
  INVX2 U8929 ( .A(n2242), .Y(n13044) );
  INVX2 U8930 ( .A(n600), .Y(n13042) );
  INVX2 U8931 ( .A(n2515), .Y(n13051) );
  INVX2 U8932 ( .A(n3062), .Y(n13049) );
  INVX2 U8933 ( .A(n3335), .Y(n13048) );
  INVX2 U8934 ( .A(n3608), .Y(n13055) );
  INVX2 U8935 ( .A(n3882), .Y(n13054) );
  INVX2 U8936 ( .A(n4155), .Y(n13053) );
  INVX2 U8937 ( .A(n4436), .Y(n13052) );
  INVX2 U8938 ( .A(n874), .Y(n13041) );
  BUFX2 U8939 ( .A(n13071), .Y(n12774) );
  BUFX2 U8940 ( .A(n13070), .Y(n12768) );
  BUFX2 U8941 ( .A(n13069), .Y(n12762) );
  BUFX2 U8942 ( .A(n13068), .Y(n12756) );
  BUFX2 U8943 ( .A(n13067), .Y(n12750) );
  BUFX2 U8944 ( .A(n13066), .Y(n12744) );
  BUFX2 U8945 ( .A(n13065), .Y(n12738) );
  BUFX2 U8946 ( .A(n13064), .Y(n12732) );
  BUFX2 U8947 ( .A(n13063), .Y(n12726) );
  BUFX2 U8948 ( .A(n13062), .Y(n12720) );
  BUFX2 U8949 ( .A(n13061), .Y(n12714) );
  BUFX2 U8950 ( .A(n13060), .Y(n12708) );
  BUFX2 U8951 ( .A(n13059), .Y(n12702) );
  BUFX2 U8952 ( .A(n13058), .Y(n12696) );
  BUFX2 U8953 ( .A(n13057), .Y(n12690) );
  BUFX2 U8954 ( .A(n13056), .Y(n12684) );
  BUFX2 U8955 ( .A(mem_access_addr[3]), .Y(n12574) );
  BUFX2 U8956 ( .A(n13071), .Y(n12775) );
  BUFX2 U8957 ( .A(n13070), .Y(n12769) );
  BUFX2 U8958 ( .A(n13069), .Y(n12763) );
  BUFX2 U8959 ( .A(n13068), .Y(n12757) );
  BUFX2 U8960 ( .A(n13067), .Y(n12751) );
  BUFX2 U8961 ( .A(n13066), .Y(n12745) );
  BUFX2 U8962 ( .A(n13065), .Y(n12739) );
  BUFX2 U8963 ( .A(n13064), .Y(n12733) );
  BUFX2 U8964 ( .A(n13063), .Y(n12727) );
  BUFX2 U8965 ( .A(n13062), .Y(n12721) );
  BUFX2 U8966 ( .A(n13061), .Y(n12715) );
  BUFX2 U8967 ( .A(n13060), .Y(n12709) );
  BUFX2 U8968 ( .A(n13059), .Y(n12703) );
  BUFX2 U8969 ( .A(n13058), .Y(n12697) );
  BUFX2 U8970 ( .A(n13057), .Y(n12691) );
  BUFX2 U8971 ( .A(n13056), .Y(n12685) );
  INVX2 U8972 ( .A(mem_access_addr[2]), .Y(n13037) );
  INVX2 U8973 ( .A(mem_access_addr[0]), .Y(n13036) );
  BUFX2 U8974 ( .A(mem_access_addr[5]), .Y(n12563) );
  BUFX2 U8975 ( .A(mem_access_addr[5]), .Y(n12562) );
  INVX2 U8976 ( .A(mem_access_addr[4]), .Y(n13038) );
  MUX2X1 U8977 ( .B(n3848), .A(n3865), .S(n12590), .Y(n3831) );
  MUX2X1 U8978 ( .B(n3900), .A(n3917), .S(n12596), .Y(n3883) );
  MUX2X1 U8979 ( .B(n3951), .A(n3968), .S(n12614), .Y(n3934) );
  MUX2X1 U8980 ( .B(n4002), .A(n4019), .S(n12601), .Y(n3985) );
  MUX2X1 U8981 ( .B(n4053), .A(n4070), .S(n12571), .Y(n4036) );
  MUX2X1 U8982 ( .B(n4104), .A(n4121), .S(n12618), .Y(n4087) );
  MUX2X1 U8983 ( .B(n4156), .A(n4175), .S(n12619), .Y(n4138) );
  MUX2X1 U8984 ( .B(n4211), .A(n4229), .S(n12603), .Y(n4193) );
  MUX2X1 U8985 ( .B(n4264), .A(n4281), .S(n12595), .Y(n4247) );
  MUX2X1 U8986 ( .B(n4316), .A(n4333), .S(n12570), .Y(n4298) );
  MUX2X1 U8987 ( .B(n4367), .A(n4385), .S(n12595), .Y(n4350) );
  MUX2X1 U8988 ( .B(n4419), .A(n8533), .S(n12619), .Y(n4402) );
  MUX2X1 U8989 ( .B(n8535), .A(n8536), .S(n12606), .Y(n8534) );
  MUX2X1 U8990 ( .B(n8538), .A(n8539), .S(n12592), .Y(n8537) );
  MUX2X1 U8991 ( .B(n8541), .A(n8542), .S(n12569), .Y(n8540) );
  MUX2X1 U8992 ( .B(n8544), .A(n8545), .S(n12614), .Y(n8543) );
  MUX2X1 U8993 ( .B(n8547), .A(n8548), .S(n12602), .Y(n8546) );
  MUX2X1 U8994 ( .B(n8550), .A(n8551), .S(n12603), .Y(n8549) );
  MUX2X1 U8995 ( .B(n8553), .A(n8554), .S(n12611), .Y(n8552) );
  MUX2X1 U8996 ( .B(n8556), .A(n8557), .S(n12572), .Y(n8555) );
  MUX2X1 U8997 ( .B(n8559), .A(n8560), .S(n12562), .Y(n8558) );
  MUX2X1 U8998 ( .B(n8562), .A(n8563), .S(n12595), .Y(n8561) );
  MUX2X1 U8999 ( .B(n8565), .A(n8566), .S(n12598), .Y(n8564) );
  MUX2X1 U9000 ( .B(n8568), .A(n8569), .S(n12617), .Y(n8567) );
  MUX2X1 U9001 ( .B(n8571), .A(n8572), .S(n12593), .Y(n8570) );
  MUX2X1 U9002 ( .B(n8574), .A(n8575), .S(n12572), .Y(n8573) );
  MUX2X1 U9003 ( .B(n8577), .A(n8578), .S(n12619), .Y(n8576) );
  MUX2X1 U9004 ( .B(n8580), .A(n8581), .S(n12620), .Y(n8579) );
  MUX2X1 U9005 ( .B(n8583), .A(n8584), .S(n12615), .Y(n8582) );
  MUX2X1 U9006 ( .B(n8586), .A(n8587), .S(n12591), .Y(n8585) );
  MUX2X1 U9007 ( .B(n8589), .A(n8590), .S(n12574), .Y(n8588) );
  MUX2X1 U9008 ( .B(n8592), .A(n8593), .S(n12601), .Y(n8591) );
  MUX2X1 U9009 ( .B(n8595), .A(n8596), .S(n12605), .Y(n8594) );
  MUX2X1 U9010 ( .B(n8598), .A(n8599), .S(n12593), .Y(n8597) );
  MUX2X1 U9011 ( .B(n8601), .A(n8602), .S(n12591), .Y(n8600) );
  MUX2X1 U9012 ( .B(n8604), .A(n8605), .S(n12569), .Y(n8603) );
  MUX2X1 U9013 ( .B(n8607), .A(n8608), .S(n12616), .Y(n8606) );
  MUX2X1 U9014 ( .B(n8610), .A(n8611), .S(n12599), .Y(n8609) );
  MUX2X1 U9015 ( .B(n8613), .A(n8614), .S(n12594), .Y(n8612) );
  MUX2X1 U9016 ( .B(n8616), .A(n8617), .S(n12614), .Y(n8615) );
  MUX2X1 U9017 ( .B(n8619), .A(n8620), .S(n12573), .Y(n8618) );
  MUX2X1 U9018 ( .B(n8622), .A(n8623), .S(n12562), .Y(n8621) );
  MUX2X1 U9019 ( .B(n8625), .A(n8626), .S(n12596), .Y(n8624) );
  MUX2X1 U9020 ( .B(n8628), .A(n8629), .S(n12618), .Y(n8627) );
  MUX2X1 U9021 ( .B(n8631), .A(n8632), .S(n12591), .Y(n8630) );
  MUX2X1 U9022 ( .B(n8634), .A(n8635), .S(n12619), .Y(n8633) );
  MUX2X1 U9023 ( .B(n8637), .A(n8638), .S(n12569), .Y(n8636) );
  MUX2X1 U9024 ( .B(n8640), .A(n8641), .S(n12591), .Y(n8639) );
  MUX2X1 U9025 ( .B(n8643), .A(n8644), .S(n12590), .Y(n8642) );
  MUX2X1 U9026 ( .B(n8646), .A(n8647), .S(n12594), .Y(n8645) );
  MUX2X1 U9027 ( .B(n8649), .A(n8650), .S(n12617), .Y(n8648) );
  MUX2X1 U9028 ( .B(n8652), .A(n8653), .S(n12571), .Y(n8651) );
  MUX2X1 U9029 ( .B(n8655), .A(n8656), .S(n12613), .Y(n8654) );
  MUX2X1 U9030 ( .B(n8658), .A(n8659), .S(n12596), .Y(n8657) );
  MUX2X1 U9031 ( .B(n8661), .A(n8662), .S(n12592), .Y(n8660) );
  MUX2X1 U9032 ( .B(n8664), .A(n8665), .S(n12615), .Y(n8663) );
  MUX2X1 U9033 ( .B(n8667), .A(n8668), .S(n12574), .Y(n8666) );
  MUX2X1 U9034 ( .B(n8670), .A(n8671), .S(n12591), .Y(n8669) );
  MUX2X1 U9035 ( .B(n8673), .A(n8674), .S(n12610), .Y(n8672) );
  MUX2X1 U9036 ( .B(n8676), .A(n8677), .S(n12595), .Y(n8675) );
  MUX2X1 U9037 ( .B(n8679), .A(n8680), .S(n12597), .Y(n8678) );
  MUX2X1 U9038 ( .B(n8682), .A(n8683), .S(n12569), .Y(n8681) );
  MUX2X1 U9039 ( .B(n8685), .A(n8686), .S(n12562), .Y(n8684) );
  MUX2X1 U9040 ( .B(n8688), .A(n8689), .S(n12597), .Y(n8687) );
  MUX2X1 U9041 ( .B(n8691), .A(n8692), .S(n12598), .Y(n8690) );
  MUX2X1 U9042 ( .B(n8694), .A(n8695), .S(n12595), .Y(n8693) );
  MUX2X1 U9043 ( .B(n8697), .A(n8698), .S(n12604), .Y(n8696) );
  MUX2X1 U9044 ( .B(n8700), .A(n8701), .S(n12574), .Y(n8699) );
  MUX2X1 U9045 ( .B(n8703), .A(n8704), .S(n12592), .Y(n8702) );
  MUX2X1 U9046 ( .B(n8706), .A(n8707), .S(n12601), .Y(n8705) );
  MUX2X1 U9047 ( .B(n8709), .A(n8710), .S(n12609), .Y(n8708) );
  MUX2X1 U9048 ( .B(n8712), .A(n8713), .S(n12614), .Y(n8711) );
  MUX2X1 U9049 ( .B(n8715), .A(n8716), .S(mem_access_addr[3]), .Y(n8714) );
  MUX2X1 U9050 ( .B(n8718), .A(n8719), .S(n12620), .Y(n8717) );
  MUX2X1 U9051 ( .B(n8721), .A(n8722), .S(n12620), .Y(n8720) );
  MUX2X1 U9052 ( .B(n8724), .A(n8725), .S(n12590), .Y(n8723) );
  MUX2X1 U9053 ( .B(n8727), .A(n8728), .S(n12606), .Y(n8726) );
  MUX2X1 U9054 ( .B(n8730), .A(n8731), .S(n12568), .Y(n8729) );
  MUX2X1 U9055 ( .B(n8733), .A(n8734), .S(n12618), .Y(n8732) );
  MUX2X1 U9056 ( .B(n8736), .A(n8737), .S(n12609), .Y(n8735) );
  MUX2X1 U9057 ( .B(n8739), .A(n8740), .S(n12612), .Y(n8738) );
  MUX2X1 U9058 ( .B(n8742), .A(n8743), .S(n12600), .Y(n8741) );
  MUX2X1 U9059 ( .B(n8745), .A(n8746), .S(n12573), .Y(n8744) );
  MUX2X1 U9060 ( .B(n8748), .A(n8749), .S(n12562), .Y(n8747) );
  MUX2X1 U9061 ( .B(n8750), .A(n8751), .S(mem_access_addr[7]), .Y(
        mem_read_data[0]) );
  MUX2X1 U9062 ( .B(n8753), .A(n8754), .S(n12613), .Y(n8752) );
  MUX2X1 U9063 ( .B(n8756), .A(n8757), .S(n12590), .Y(n8755) );
  MUX2X1 U9064 ( .B(n8759), .A(n8760), .S(n12617), .Y(n8758) );
  MUX2X1 U9065 ( .B(n8762), .A(n8763), .S(n12607), .Y(n8761) );
  MUX2X1 U9066 ( .B(n8765), .A(n8766), .S(n12571), .Y(n8764) );
  MUX2X1 U9067 ( .B(n8768), .A(n8769), .S(n12606), .Y(n8767) );
  MUX2X1 U9068 ( .B(n8771), .A(n8772), .S(n12592), .Y(n8770) );
  MUX2X1 U9069 ( .B(n8774), .A(n8775), .S(n12604), .Y(n8773) );
  MUX2X1 U9070 ( .B(n8777), .A(n8778), .S(n12619), .Y(n8776) );
  MUX2X1 U9071 ( .B(n8780), .A(n8781), .S(mem_access_addr[3]), .Y(n8779) );
  MUX2X1 U9072 ( .B(n8783), .A(n8784), .S(n12607), .Y(n8782) );
  MUX2X1 U9073 ( .B(n8786), .A(n8787), .S(n12608), .Y(n8785) );
  MUX2X1 U9074 ( .B(n8789), .A(n8790), .S(n12591), .Y(n8788) );
  MUX2X1 U9075 ( .B(n8792), .A(n8793), .S(n12590), .Y(n8791) );
  MUX2X1 U9076 ( .B(n8795), .A(n8796), .S(n12570), .Y(n8794) );
  MUX2X1 U9077 ( .B(n8798), .A(n8799), .S(n12612), .Y(n8797) );
  MUX2X1 U9078 ( .B(n8801), .A(n8802), .S(n12612), .Y(n8800) );
  MUX2X1 U9079 ( .B(n8804), .A(n8805), .S(n12617), .Y(n8803) );
  MUX2X1 U9080 ( .B(n8807), .A(n8808), .S(n12612), .Y(n8806) );
  MUX2X1 U9081 ( .B(n8810), .A(n8811), .S(n12568), .Y(n8809) );
  MUX2X1 U9082 ( .B(n8813), .A(n8814), .S(n12563), .Y(n8812) );
  MUX2X1 U9083 ( .B(n8816), .A(n8817), .S(n12596), .Y(n8815) );
  MUX2X1 U9084 ( .B(n8819), .A(n8820), .S(n12605), .Y(n8818) );
  MUX2X1 U9085 ( .B(n8822), .A(n8823), .S(n12619), .Y(n8821) );
  MUX2X1 U9086 ( .B(n8825), .A(n8826), .S(n12601), .Y(n8824) );
  MUX2X1 U9087 ( .B(n8828), .A(n8829), .S(n12570), .Y(n8827) );
  MUX2X1 U9088 ( .B(n8831), .A(n8832), .S(mem_access_addr[1]), .Y(n8830) );
  MUX2X1 U9089 ( .B(n8834), .A(n8835), .S(n12616), .Y(n8833) );
  MUX2X1 U9090 ( .B(n8837), .A(n8838), .S(n12606), .Y(n8836) );
  MUX2X1 U9091 ( .B(n8840), .A(n8841), .S(n12604), .Y(n8839) );
  MUX2X1 U9092 ( .B(n8843), .A(n8844), .S(mem_access_addr[3]), .Y(n8842) );
  MUX2X1 U9093 ( .B(n8846), .A(n8847), .S(n12596), .Y(n8845) );
  MUX2X1 U9094 ( .B(n8849), .A(n8850), .S(mem_access_addr[1]), .Y(n8848) );
  MUX2X1 U9095 ( .B(n8852), .A(n8853), .S(n12597), .Y(n8851) );
  MUX2X1 U9096 ( .B(n8855), .A(n8856), .S(n12601), .Y(n8854) );
  MUX2X1 U9097 ( .B(n8858), .A(n8859), .S(n12570), .Y(n8857) );
  MUX2X1 U9098 ( .B(n8861), .A(n8862), .S(mem_access_addr[1]), .Y(n8860) );
  MUX2X1 U9099 ( .B(n8864), .A(n8865), .S(n12603), .Y(n8863) );
  MUX2X1 U9100 ( .B(n8867), .A(n8868), .S(n12615), .Y(n8866) );
  MUX2X1 U9101 ( .B(n8870), .A(n8871), .S(n12609), .Y(n8869) );
  MUX2X1 U9102 ( .B(n8873), .A(n8874), .S(n12570), .Y(n8872) );
  MUX2X1 U9103 ( .B(n8876), .A(n8877), .S(n12563), .Y(n8875) );
  MUX2X1 U9104 ( .B(n8879), .A(n8880), .S(n12594), .Y(n8878) );
  MUX2X1 U9105 ( .B(n8882), .A(n8883), .S(n12608), .Y(n8881) );
  MUX2X1 U9106 ( .B(n8885), .A(n8886), .S(n12594), .Y(n8884) );
  MUX2X1 U9107 ( .B(n8888), .A(n8889), .S(n12594), .Y(n8887) );
  MUX2X1 U9108 ( .B(n8891), .A(n8892), .S(n12574), .Y(n8890) );
  MUX2X1 U9109 ( .B(n8894), .A(n8895), .S(n12605), .Y(n8893) );
  MUX2X1 U9110 ( .B(n8897), .A(n8898), .S(n12607), .Y(n8896) );
  MUX2X1 U9111 ( .B(n8900), .A(n8901), .S(n12600), .Y(n8899) );
  MUX2X1 U9112 ( .B(n8903), .A(n8904), .S(n12591), .Y(n8902) );
  MUX2X1 U9113 ( .B(n8906), .A(n8907), .S(n12573), .Y(n8905) );
  MUX2X1 U9114 ( .B(n8909), .A(n8910), .S(n12615), .Y(n8908) );
  MUX2X1 U9115 ( .B(n8912), .A(n8913), .S(n12608), .Y(n8911) );
  MUX2X1 U9116 ( .B(n8915), .A(n8916), .S(n12613), .Y(n8914) );
  MUX2X1 U9117 ( .B(n8918), .A(n8919), .S(n12617), .Y(n8917) );
  MUX2X1 U9118 ( .B(n8921), .A(n8922), .S(n12570), .Y(n8920) );
  MUX2X1 U9119 ( .B(n8924), .A(n8925), .S(n12603), .Y(n8923) );
  MUX2X1 U9120 ( .B(n8927), .A(n8928), .S(n12603), .Y(n8926) );
  MUX2X1 U9121 ( .B(n8930), .A(n8931), .S(n12604), .Y(n8929) );
  MUX2X1 U9122 ( .B(n8933), .A(n8934), .S(n12599), .Y(n8932) );
  MUX2X1 U9123 ( .B(n8936), .A(n8937), .S(n12570), .Y(n8935) );
  MUX2X1 U9124 ( .B(n8939), .A(n8940), .S(n12563), .Y(n8938) );
  MUX2X1 U9125 ( .B(n8942), .A(n8943), .S(n12612), .Y(n8941) );
  MUX2X1 U9126 ( .B(n8945), .A(n8946), .S(n12613), .Y(n8944) );
  MUX2X1 U9127 ( .B(n8948), .A(n8949), .S(n12605), .Y(n8947) );
  MUX2X1 U9128 ( .B(n8951), .A(n8952), .S(n12610), .Y(n8950) );
  MUX2X1 U9129 ( .B(n8954), .A(n8955), .S(n12574), .Y(n8953) );
  MUX2X1 U9130 ( .B(n8957), .A(n8958), .S(n12599), .Y(n8956) );
  MUX2X1 U9131 ( .B(n8960), .A(n8961), .S(n12597), .Y(n8959) );
  MUX2X1 U9132 ( .B(n8963), .A(n8964), .S(n12620), .Y(n8962) );
  MUX2X1 U9133 ( .B(n8966), .A(n8967), .S(n12604), .Y(n8965) );
  MUX2X1 U9134 ( .B(n8969), .A(n8970), .S(n12569), .Y(n8968) );
  MUX2X1 U9135 ( .B(n8972), .A(n8973), .S(n12613), .Y(n8971) );
  MUX2X1 U9136 ( .B(n8975), .A(n8976), .S(n12616), .Y(n8974) );
  MUX2X1 U9137 ( .B(n8978), .A(n8979), .S(n12595), .Y(n8977) );
  MUX2X1 U9138 ( .B(n8981), .A(n8982), .S(n12602), .Y(n8980) );
  MUX2X1 U9139 ( .B(n8984), .A(n8985), .S(n12574), .Y(n8983) );
  MUX2X1 U9140 ( .B(n8987), .A(n8988), .S(n12618), .Y(n8986) );
  MUX2X1 U9141 ( .B(n8990), .A(n8991), .S(n12607), .Y(n8989) );
  MUX2X1 U9142 ( .B(n8993), .A(n8994), .S(n12598), .Y(n8992) );
  MUX2X1 U9143 ( .B(n8996), .A(n8997), .S(n12590), .Y(n8995) );
  MUX2X1 U9144 ( .B(n8999), .A(n9000), .S(n12574), .Y(n8998) );
  MUX2X1 U9145 ( .B(n9002), .A(n9003), .S(n12563), .Y(n9001) );
  MUX2X1 U9146 ( .B(n9004), .A(n9005), .S(mem_access_addr[7]), .Y(
        mem_read_data[1]) );
  MUX2X1 U9147 ( .B(n9007), .A(n9008), .S(n12598), .Y(n9006) );
  MUX2X1 U9148 ( .B(n9010), .A(n9011), .S(n12597), .Y(n9009) );
  MUX2X1 U9149 ( .B(n9013), .A(n9014), .S(n12611), .Y(n9012) );
  MUX2X1 U9150 ( .B(n9016), .A(n9017), .S(n12610), .Y(n9015) );
  MUX2X1 U9151 ( .B(n9019), .A(n9020), .S(n12570), .Y(n9018) );
  MUX2X1 U9152 ( .B(n9022), .A(n9023), .S(n12606), .Y(n9021) );
  MUX2X1 U9153 ( .B(n9025), .A(n9026), .S(n12598), .Y(n9024) );
  MUX2X1 U9154 ( .B(n9028), .A(n9029), .S(n12613), .Y(n9027) );
  MUX2X1 U9155 ( .B(n9031), .A(n9032), .S(n12615), .Y(n9030) );
  MUX2X1 U9156 ( .B(n9034), .A(n9035), .S(n12574), .Y(n9033) );
  MUX2X1 U9157 ( .B(n9037), .A(n9038), .S(n12594), .Y(n9036) );
  MUX2X1 U9158 ( .B(n9040), .A(n9041), .S(n12599), .Y(n9039) );
  MUX2X1 U9159 ( .B(n9043), .A(n9044), .S(n12592), .Y(n9042) );
  MUX2X1 U9160 ( .B(n9046), .A(n9047), .S(n12608), .Y(n9045) );
  MUX2X1 U9161 ( .B(n9049), .A(n9050), .S(n12574), .Y(n9048) );
  MUX2X1 U9162 ( .B(n9052), .A(n9053), .S(n12615), .Y(n9051) );
  MUX2X1 U9163 ( .B(n9055), .A(n9056), .S(n12600), .Y(n9054) );
  MUX2X1 U9164 ( .B(n9058), .A(n9059), .S(n12613), .Y(n9057) );
  MUX2X1 U9165 ( .B(n9061), .A(n9062), .S(n12595), .Y(n9060) );
  MUX2X1 U9166 ( .B(n9064), .A(n9065), .S(n12574), .Y(n9063) );
  MUX2X1 U9167 ( .B(n9067), .A(n9068), .S(n12563), .Y(n9066) );
  MUX2X1 U9168 ( .B(n9070), .A(n9071), .S(n12607), .Y(n9069) );
  MUX2X1 U9169 ( .B(n9073), .A(n9074), .S(n12613), .Y(n9072) );
  MUX2X1 U9170 ( .B(n9076), .A(n9077), .S(n12607), .Y(n9075) );
  MUX2X1 U9171 ( .B(n9079), .A(n9080), .S(n12606), .Y(n9078) );
  MUX2X1 U9172 ( .B(n9082), .A(n9083), .S(n12574), .Y(n9081) );
  MUX2X1 U9173 ( .B(n9085), .A(n9086), .S(n12619), .Y(n9084) );
  MUX2X1 U9174 ( .B(n9088), .A(n9089), .S(n12598), .Y(n9087) );
  MUX2X1 U9175 ( .B(n9091), .A(n9092), .S(n12602), .Y(n9090) );
  MUX2X1 U9176 ( .B(n9094), .A(n9095), .S(n12607), .Y(n9093) );
  MUX2X1 U9177 ( .B(n9097), .A(n9098), .S(mem_access_addr[3]), .Y(n9096) );
  MUX2X1 U9178 ( .B(n9100), .A(n9101), .S(n12604), .Y(n9099) );
  MUX2X1 U9179 ( .B(n9103), .A(n9104), .S(mem_access_addr[1]), .Y(n9102) );
  MUX2X1 U9180 ( .B(n9106), .A(n9107), .S(n12594), .Y(n9105) );
  MUX2X1 U9181 ( .B(n9109), .A(n9110), .S(n12619), .Y(n9108) );
  MUX2X1 U9182 ( .B(n9112), .A(n9113), .S(n12570), .Y(n9111) );
  MUX2X1 U9183 ( .B(n9115), .A(n9116), .S(n12618), .Y(n9114) );
  MUX2X1 U9184 ( .B(n9118), .A(n9119), .S(n12595), .Y(n9117) );
  MUX2X1 U9185 ( .B(n9121), .A(n9122), .S(n12608), .Y(n9120) );
  MUX2X1 U9186 ( .B(n9124), .A(n9125), .S(n12593), .Y(n9123) );
  MUX2X1 U9187 ( .B(n9127), .A(n9128), .S(n12574), .Y(n9126) );
  MUX2X1 U9188 ( .B(n9130), .A(n9131), .S(n12563), .Y(n9129) );
  MUX2X1 U9189 ( .B(n9133), .A(n9134), .S(n12605), .Y(n9132) );
  MUX2X1 U9190 ( .B(n9136), .A(n9137), .S(n12609), .Y(n9135) );
  MUX2X1 U9191 ( .B(n9139), .A(n9140), .S(n12590), .Y(n9138) );
  MUX2X1 U9192 ( .B(n9142), .A(n9143), .S(n12605), .Y(n9141) );
  MUX2X1 U9193 ( .B(n9145), .A(n9146), .S(n12568), .Y(n9144) );
  MUX2X1 U9194 ( .B(n9148), .A(n9149), .S(n12602), .Y(n9147) );
  MUX2X1 U9195 ( .B(n9151), .A(n9152), .S(n12614), .Y(n9150) );
  MUX2X1 U9196 ( .B(n9154), .A(n9155), .S(n12600), .Y(n9153) );
  MUX2X1 U9197 ( .B(n9157), .A(n9158), .S(n12609), .Y(n9156) );
  MUX2X1 U9198 ( .B(n9160), .A(n9161), .S(n12568), .Y(n9159) );
  MUX2X1 U9199 ( .B(n9163), .A(n9164), .S(n12614), .Y(n9162) );
  MUX2X1 U9200 ( .B(n9166), .A(n9167), .S(n12604), .Y(n9165) );
  MUX2X1 U9201 ( .B(n9169), .A(n9170), .S(n12592), .Y(n9168) );
  MUX2X1 U9202 ( .B(n9172), .A(n9173), .S(n12591), .Y(n9171) );
  MUX2X1 U9203 ( .B(n9175), .A(n9176), .S(n12568), .Y(n9174) );
  MUX2X1 U9204 ( .B(n9178), .A(n9179), .S(n12591), .Y(n9177) );
  MUX2X1 U9205 ( .B(n9181), .A(n9182), .S(n12606), .Y(n9180) );
  MUX2X1 U9206 ( .B(n9184), .A(n9185), .S(n12599), .Y(n9183) );
  MUX2X1 U9207 ( .B(n9187), .A(n9188), .S(n12616), .Y(n9186) );
  MUX2X1 U9208 ( .B(n9190), .A(n9191), .S(n12568), .Y(n9189) );
  MUX2X1 U9209 ( .B(n9193), .A(n9194), .S(n12563), .Y(n9192) );
  MUX2X1 U9210 ( .B(n9196), .A(n9197), .S(n12609), .Y(n9195) );
  MUX2X1 U9211 ( .B(n9199), .A(n9200), .S(n12591), .Y(n9198) );
  MUX2X1 U9212 ( .B(n9202), .A(n9203), .S(n12593), .Y(n9201) );
  MUX2X1 U9213 ( .B(n9205), .A(n9206), .S(n12620), .Y(n9204) );
  MUX2X1 U9214 ( .B(n9208), .A(n9209), .S(n12568), .Y(n9207) );
  MUX2X1 U9215 ( .B(n9211), .A(n9212), .S(n12618), .Y(n9210) );
  MUX2X1 U9216 ( .B(n9214), .A(n9215), .S(n12620), .Y(n9213) );
  MUX2X1 U9217 ( .B(n9217), .A(n9218), .S(n12618), .Y(n9216) );
  MUX2X1 U9218 ( .B(n9220), .A(n9221), .S(n12593), .Y(n9219) );
  MUX2X1 U9219 ( .B(n9223), .A(n9224), .S(n12571), .Y(n9222) );
  MUX2X1 U9220 ( .B(n9226), .A(n9227), .S(n12604), .Y(n9225) );
  MUX2X1 U9221 ( .B(n9229), .A(n9230), .S(n12615), .Y(n9228) );
  MUX2X1 U9222 ( .B(n9232), .A(n9233), .S(n12593), .Y(n9231) );
  MUX2X1 U9223 ( .B(n9235), .A(n9236), .S(n12614), .Y(n9234) );
  MUX2X1 U9224 ( .B(n9238), .A(n9239), .S(n12568), .Y(n9237) );
  MUX2X1 U9225 ( .B(n9241), .A(n9242), .S(n12599), .Y(n9240) );
  MUX2X1 U9226 ( .B(n9244), .A(n9245), .S(n12606), .Y(n9243) );
  MUX2X1 U9227 ( .B(n9247), .A(n9248), .S(n12604), .Y(n9246) );
  MUX2X1 U9228 ( .B(n9250), .A(n9251), .S(n12610), .Y(n9249) );
  MUX2X1 U9229 ( .B(n9253), .A(n9254), .S(n12568), .Y(n9252) );
  MUX2X1 U9230 ( .B(n9256), .A(n9257), .S(n12563), .Y(n9255) );
  MUX2X1 U9231 ( .B(n9258), .A(n9259), .S(mem_access_addr[7]), .Y(
        mem_read_data[2]) );
  MUX2X1 U9232 ( .B(n9261), .A(n9262), .S(n12596), .Y(n9260) );
  MUX2X1 U9233 ( .B(n9264), .A(n9265), .S(n12600), .Y(n9263) );
  MUX2X1 U9234 ( .B(n9267), .A(n9268), .S(n12613), .Y(n9266) );
  MUX2X1 U9235 ( .B(n9270), .A(n9271), .S(n12590), .Y(n9269) );
  MUX2X1 U9236 ( .B(n9273), .A(n9274), .S(n12568), .Y(n9272) );
  MUX2X1 U9237 ( .B(n9276), .A(n9277), .S(n12597), .Y(n9275) );
  MUX2X1 U9238 ( .B(n9279), .A(n9280), .S(n12596), .Y(n9278) );
  MUX2X1 U9239 ( .B(n9282), .A(n9283), .S(n12594), .Y(n9281) );
  MUX2X1 U9240 ( .B(n9285), .A(n9286), .S(n12605), .Y(n9284) );
  MUX2X1 U9241 ( .B(n9288), .A(n9289), .S(n12573), .Y(n9287) );
  MUX2X1 U9242 ( .B(n9291), .A(n9292), .S(n12605), .Y(n9290) );
  MUX2X1 U9243 ( .B(n9294), .A(n9295), .S(n12619), .Y(n9293) );
  MUX2X1 U9244 ( .B(n9297), .A(n9298), .S(n12596), .Y(n9296) );
  MUX2X1 U9245 ( .B(n9300), .A(n9301), .S(n12607), .Y(n9299) );
  MUX2X1 U9246 ( .B(n9303), .A(n9304), .S(n12568), .Y(n9302) );
  MUX2X1 U9247 ( .B(n9306), .A(n9307), .S(n12610), .Y(n9305) );
  MUX2X1 U9248 ( .B(n9309), .A(n9310), .S(n12606), .Y(n9308) );
  MUX2X1 U9249 ( .B(n9312), .A(n9313), .S(n12601), .Y(n9311) );
  MUX2X1 U9250 ( .B(n9315), .A(n9316), .S(n12603), .Y(n9314) );
  MUX2X1 U9251 ( .B(n9318), .A(n9319), .S(n12568), .Y(n9317) );
  MUX2X1 U9252 ( .B(n9321), .A(n9322), .S(n12563), .Y(n9320) );
  MUX2X1 U9253 ( .B(n9324), .A(n9325), .S(n12598), .Y(n9323) );
  MUX2X1 U9254 ( .B(n9327), .A(n9328), .S(n12620), .Y(n9326) );
  MUX2X1 U9255 ( .B(n9330), .A(n9331), .S(n12619), .Y(n9329) );
  MUX2X1 U9256 ( .B(n9333), .A(n9334), .S(n12590), .Y(n9332) );
  MUX2X1 U9257 ( .B(n9336), .A(n9337), .S(n12574), .Y(n9335) );
  MUX2X1 U9258 ( .B(n9339), .A(n9340), .S(n12615), .Y(n9338) );
  MUX2X1 U9259 ( .B(n9342), .A(n9343), .S(n12611), .Y(n9341) );
  MUX2X1 U9260 ( .B(n9345), .A(n9346), .S(n12618), .Y(n9344) );
  MUX2X1 U9261 ( .B(n9348), .A(n9349), .S(n12620), .Y(n9347) );
  MUX2X1 U9262 ( .B(n9351), .A(n9352), .S(n12571), .Y(n9350) );
  MUX2X1 U9263 ( .B(n9354), .A(n9355), .S(n12591), .Y(n9353) );
  MUX2X1 U9264 ( .B(n9357), .A(n9358), .S(n12618), .Y(n9356) );
  MUX2X1 U9265 ( .B(n9360), .A(n9361), .S(n12595), .Y(n9359) );
  MUX2X1 U9266 ( .B(n9363), .A(n9364), .S(n12603), .Y(n9362) );
  MUX2X1 U9267 ( .B(n9366), .A(n9367), .S(n12571), .Y(n9365) );
  MUX2X1 U9268 ( .B(n9369), .A(n9370), .S(mem_access_addr[1]), .Y(n9368) );
  MUX2X1 U9269 ( .B(n9372), .A(n9373), .S(n12594), .Y(n9371) );
  MUX2X1 U9270 ( .B(n9375), .A(n9376), .S(n12605), .Y(n9374) );
  MUX2X1 U9271 ( .B(n9378), .A(n9379), .S(n12620), .Y(n9377) );
  MUX2X1 U9272 ( .B(n9381), .A(n9382), .S(n12572), .Y(n9380) );
  MUX2X1 U9273 ( .B(n9384), .A(n9385), .S(n12563), .Y(n9383) );
  MUX2X1 U9274 ( .B(n9387), .A(n9388), .S(n12598), .Y(n9386) );
  MUX2X1 U9275 ( .B(n9390), .A(n9391), .S(n12592), .Y(n9389) );
  MUX2X1 U9276 ( .B(n9393), .A(n9394), .S(n12591), .Y(n9392) );
  MUX2X1 U9277 ( .B(n9396), .A(n9397), .S(n12610), .Y(n9395) );
  MUX2X1 U9278 ( .B(n9399), .A(n9400), .S(n12571), .Y(n9398) );
  MUX2X1 U9279 ( .B(n9402), .A(n9403), .S(n12620), .Y(n9401) );
  MUX2X1 U9280 ( .B(n9405), .A(n9406), .S(n12607), .Y(n9404) );
  MUX2X1 U9281 ( .B(n9408), .A(n9409), .S(n12598), .Y(n9407) );
  MUX2X1 U9282 ( .B(n9411), .A(n9412), .S(n12611), .Y(n9410) );
  MUX2X1 U9283 ( .B(n9414), .A(n9415), .S(n12571), .Y(n9413) );
  MUX2X1 U9284 ( .B(n9417), .A(n9418), .S(n12606), .Y(n9416) );
  MUX2X1 U9285 ( .B(n9420), .A(n9421), .S(n12616), .Y(n9419) );
  MUX2X1 U9286 ( .B(n9423), .A(n9424), .S(n12591), .Y(n9422) );
  MUX2X1 U9287 ( .B(n9426), .A(n9427), .S(n12600), .Y(n9425) );
  MUX2X1 U9288 ( .B(n9429), .A(n9430), .S(n12568), .Y(n9428) );
  MUX2X1 U9289 ( .B(n9432), .A(n9433), .S(n12612), .Y(n9431) );
  MUX2X1 U9290 ( .B(n9435), .A(n9436), .S(n12605), .Y(n9434) );
  MUX2X1 U9291 ( .B(n9438), .A(n9439), .S(n12591), .Y(n9437) );
  MUX2X1 U9292 ( .B(n9441), .A(n9442), .S(n12597), .Y(n9440) );
  MUX2X1 U9293 ( .B(n9444), .A(n9445), .S(n12568), .Y(n9443) );
  MUX2X1 U9294 ( .B(n9447), .A(n9448), .S(n12563), .Y(n9446) );
  MUX2X1 U9295 ( .B(n9450), .A(n9451), .S(n12620), .Y(n9449) );
  MUX2X1 U9296 ( .B(n9453), .A(n9454), .S(n12592), .Y(n9452) );
  MUX2X1 U9297 ( .B(n9456), .A(n9457), .S(n12610), .Y(n9455) );
  MUX2X1 U9298 ( .B(n9459), .A(n9460), .S(n12593), .Y(n9458) );
  MUX2X1 U9299 ( .B(n9462), .A(n9463), .S(mem_access_addr[3]), .Y(n9461) );
  MUX2X1 U9300 ( .B(n9465), .A(n9466), .S(n12614), .Y(n9464) );
  MUX2X1 U9301 ( .B(n9468), .A(n9469), .S(n12618), .Y(n9467) );
  MUX2X1 U9302 ( .B(n9471), .A(n9472), .S(n12592), .Y(n9470) );
  MUX2X1 U9303 ( .B(n9474), .A(n9475), .S(n12599), .Y(n9473) );
  MUX2X1 U9304 ( .B(n9477), .A(n9478), .S(n12573), .Y(n9476) );
  MUX2X1 U9305 ( .B(n9480), .A(n9481), .S(n12590), .Y(n9479) );
  MUX2X1 U9306 ( .B(n9483), .A(n9484), .S(n12617), .Y(n9482) );
  MUX2X1 U9307 ( .B(n9486), .A(n9487), .S(n12590), .Y(n9485) );
  MUX2X1 U9308 ( .B(n9489), .A(n9490), .S(n12593), .Y(n9488) );
  MUX2X1 U9309 ( .B(n9492), .A(n9493), .S(n12569), .Y(n9491) );
  MUX2X1 U9310 ( .B(n9495), .A(n9496), .S(n12619), .Y(n9494) );
  MUX2X1 U9311 ( .B(n9498), .A(n9499), .S(n12607), .Y(n9497) );
  MUX2X1 U9312 ( .B(n9501), .A(n9502), .S(n12592), .Y(n9500) );
  MUX2X1 U9313 ( .B(n9504), .A(n9505), .S(n12600), .Y(n9503) );
  MUX2X1 U9314 ( .B(n9507), .A(n9508), .S(n12571), .Y(n9506) );
  MUX2X1 U9315 ( .B(n9510), .A(n9511), .S(n12563), .Y(n9509) );
  MUX2X1 U9316 ( .B(n9512), .A(n9513), .S(mem_access_addr[7]), .Y(
        mem_read_data[3]) );
  MUX2X1 U9317 ( .B(n9515), .A(n9516), .S(n12602), .Y(n9514) );
  MUX2X1 U9318 ( .B(n9518), .A(n9519), .S(n12593), .Y(n9517) );
  MUX2X1 U9319 ( .B(n9521), .A(n9522), .S(n12604), .Y(n9520) );
  MUX2X1 U9320 ( .B(n9524), .A(n9525), .S(n12601), .Y(n9523) );
  MUX2X1 U9321 ( .B(n9527), .A(n9528), .S(n12573), .Y(n9526) );
  MUX2X1 U9322 ( .B(n9530), .A(n9531), .S(n12611), .Y(n9529) );
  MUX2X1 U9323 ( .B(n9533), .A(n9534), .S(n12618), .Y(n9532) );
  MUX2X1 U9324 ( .B(n9536), .A(n9537), .S(n12612), .Y(n9535) );
  MUX2X1 U9325 ( .B(n9539), .A(n9540), .S(mem_access_addr[1]), .Y(n9538) );
  MUX2X1 U9326 ( .B(n9542), .A(n9543), .S(n12573), .Y(n9541) );
  MUX2X1 U9327 ( .B(n9545), .A(n9546), .S(n12620), .Y(n9544) );
  MUX2X1 U9328 ( .B(n9548), .A(n9549), .S(n12612), .Y(n9547) );
  MUX2X1 U9329 ( .B(n9551), .A(n9552), .S(n12614), .Y(n9550) );
  MUX2X1 U9330 ( .B(n9554), .A(n9555), .S(n12611), .Y(n9553) );
  MUX2X1 U9331 ( .B(n9557), .A(n9558), .S(n12568), .Y(n9556) );
  MUX2X1 U9332 ( .B(n9560), .A(n9561), .S(n12596), .Y(n9559) );
  MUX2X1 U9333 ( .B(n9563), .A(n9564), .S(n12592), .Y(n9562) );
  MUX2X1 U9334 ( .B(n9566), .A(n9567), .S(n12617), .Y(n9565) );
  MUX2X1 U9335 ( .B(n9569), .A(n9570), .S(n12594), .Y(n9568) );
  MUX2X1 U9336 ( .B(n9572), .A(n9573), .S(n12569), .Y(n9571) );
  MUX2X1 U9337 ( .B(n9575), .A(n9576), .S(n12562), .Y(n9574) );
  MUX2X1 U9338 ( .B(n9578), .A(n9579), .S(n12602), .Y(n9577) );
  MUX2X1 U9339 ( .B(n9581), .A(n9582), .S(n12608), .Y(n9580) );
  MUX2X1 U9340 ( .B(n9584), .A(n9585), .S(n12595), .Y(n9583) );
  MUX2X1 U9341 ( .B(n9587), .A(n9588), .S(n12614), .Y(n9586) );
  MUX2X1 U9342 ( .B(n9590), .A(n9591), .S(mem_access_addr[3]), .Y(n9589) );
  MUX2X1 U9343 ( .B(n9593), .A(n9594), .S(n12616), .Y(n9592) );
  MUX2X1 U9344 ( .B(n9596), .A(n9597), .S(n12611), .Y(n9595) );
  MUX2X1 U9345 ( .B(n9599), .A(n9600), .S(n12609), .Y(n9598) );
  MUX2X1 U9346 ( .B(n9602), .A(n9603), .S(n12618), .Y(n9601) );
  MUX2X1 U9347 ( .B(n9605), .A(n9606), .S(n12569), .Y(n9604) );
  MUX2X1 U9348 ( .B(n9608), .A(n9609), .S(n12601), .Y(n9607) );
  MUX2X1 U9349 ( .B(n9611), .A(n9612), .S(n12599), .Y(n9610) );
  MUX2X1 U9350 ( .B(n9614), .A(n9615), .S(n12597), .Y(n9613) );
  MUX2X1 U9351 ( .B(n9617), .A(n9618), .S(n12617), .Y(n9616) );
  MUX2X1 U9352 ( .B(n9620), .A(n9621), .S(n12568), .Y(n9619) );
  MUX2X1 U9353 ( .B(n9623), .A(n9624), .S(n12620), .Y(n9622) );
  MUX2X1 U9354 ( .B(n9626), .A(n9627), .S(n12617), .Y(n9625) );
  MUX2X1 U9355 ( .B(n9629), .A(n9630), .S(n12592), .Y(n9628) );
  MUX2X1 U9356 ( .B(n9632), .A(n9633), .S(n12595), .Y(n9631) );
  MUX2X1 U9357 ( .B(n9635), .A(n9636), .S(n12569), .Y(n9634) );
  MUX2X1 U9358 ( .B(n9638), .A(n9639), .S(n12562), .Y(n9637) );
  MUX2X1 U9359 ( .B(n9641), .A(n9642), .S(n12615), .Y(n9640) );
  MUX2X1 U9360 ( .B(n9644), .A(n9645), .S(n12611), .Y(n9643) );
  MUX2X1 U9361 ( .B(n9647), .A(n9648), .S(n12602), .Y(n9646) );
  MUX2X1 U9362 ( .B(n9650), .A(n9651), .S(n12612), .Y(n9649) );
  MUX2X1 U9363 ( .B(n9653), .A(n9654), .S(n12572), .Y(n9652) );
  MUX2X1 U9364 ( .B(n9656), .A(n9657), .S(n12613), .Y(n9655) );
  MUX2X1 U9365 ( .B(n9659), .A(n9660), .S(n12594), .Y(n9658) );
  MUX2X1 U9366 ( .B(n9662), .A(n9663), .S(n12602), .Y(n9661) );
  MUX2X1 U9367 ( .B(n9665), .A(n9666), .S(n12603), .Y(n9664) );
  MUX2X1 U9368 ( .B(n9668), .A(n9669), .S(n12570), .Y(n9667) );
  MUX2X1 U9369 ( .B(n9671), .A(n9672), .S(n12608), .Y(n9670) );
  MUX2X1 U9370 ( .B(n9674), .A(n9675), .S(n12610), .Y(n9673) );
  MUX2X1 U9371 ( .B(n9677), .A(n9678), .S(n12604), .Y(n9676) );
  MUX2X1 U9372 ( .B(n9680), .A(n9681), .S(n12607), .Y(n9679) );
  MUX2X1 U9373 ( .B(n9683), .A(n9684), .S(n12571), .Y(n9682) );
  MUX2X1 U9374 ( .B(n9686), .A(n9687), .S(n12607), .Y(n9685) );
  MUX2X1 U9375 ( .B(n9689), .A(n9690), .S(n12598), .Y(n9688) );
  MUX2X1 U9376 ( .B(n9692), .A(n9693), .S(n12594), .Y(n9691) );
  MUX2X1 U9377 ( .B(n9695), .A(n9696), .S(n12593), .Y(n9694) );
  MUX2X1 U9378 ( .B(n9698), .A(n9699), .S(n12572), .Y(n9697) );
  MUX2X1 U9379 ( .B(n9701), .A(n9702), .S(n12562), .Y(n9700) );
  MUX2X1 U9380 ( .B(n9704), .A(n9705), .S(n12611), .Y(n9703) );
  MUX2X1 U9381 ( .B(n9707), .A(n9708), .S(n12605), .Y(n9706) );
  MUX2X1 U9382 ( .B(n9710), .A(n9711), .S(n12597), .Y(n9709) );
  MUX2X1 U9383 ( .B(n9713), .A(n9714), .S(n12617), .Y(n9712) );
  MUX2X1 U9384 ( .B(n9716), .A(n9717), .S(mem_access_addr[3]), .Y(n9715) );
  MUX2X1 U9385 ( .B(n9719), .A(n9720), .S(n12594), .Y(n9718) );
  MUX2X1 U9386 ( .B(n9722), .A(n9723), .S(n12601), .Y(n9721) );
  MUX2X1 U9387 ( .B(n9725), .A(n9726), .S(n12607), .Y(n9724) );
  MUX2X1 U9388 ( .B(n9728), .A(n9729), .S(n12619), .Y(n9727) );
  MUX2X1 U9389 ( .B(n9731), .A(n9732), .S(n12571), .Y(n9730) );
  MUX2X1 U9390 ( .B(n9734), .A(n9735), .S(n12609), .Y(n9733) );
  MUX2X1 U9391 ( .B(n9737), .A(n9738), .S(n12593), .Y(n9736) );
  MUX2X1 U9392 ( .B(n9740), .A(n9741), .S(n12593), .Y(n9739) );
  MUX2X1 U9393 ( .B(n9743), .A(n9744), .S(n12617), .Y(n9742) );
  MUX2X1 U9394 ( .B(n9746), .A(n9747), .S(n12569), .Y(n9745) );
  MUX2X1 U9395 ( .B(n9749), .A(n9750), .S(n12601), .Y(n9748) );
  MUX2X1 U9396 ( .B(n9752), .A(n9753), .S(n12618), .Y(n9751) );
  MUX2X1 U9397 ( .B(n9755), .A(n9756), .S(n12599), .Y(n9754) );
  MUX2X1 U9398 ( .B(n9758), .A(n9759), .S(n12597), .Y(n9757) );
  MUX2X1 U9399 ( .B(n9761), .A(n9762), .S(mem_access_addr[3]), .Y(n9760) );
  MUX2X1 U9400 ( .B(n9764), .A(n9765), .S(n12562), .Y(n9763) );
  MUX2X1 U9401 ( .B(n9766), .A(n9767), .S(mem_access_addr[7]), .Y(
        mem_read_data[4]) );
  MUX2X1 U9402 ( .B(n9769), .A(n9770), .S(n12595), .Y(n9768) );
  MUX2X1 U9403 ( .B(n9772), .A(n9773), .S(n12612), .Y(n9771) );
  MUX2X1 U9404 ( .B(n9775), .A(n9776), .S(n12590), .Y(n9774) );
  MUX2X1 U9405 ( .B(n9778), .A(n9779), .S(n12616), .Y(n9777) );
  MUX2X1 U9406 ( .B(n9781), .A(n9782), .S(n12571), .Y(n9780) );
  MUX2X1 U9407 ( .B(n9784), .A(n9785), .S(n12590), .Y(n9783) );
  MUX2X1 U9408 ( .B(n9787), .A(n9788), .S(n12600), .Y(n9786) );
  MUX2X1 U9409 ( .B(n9790), .A(n9791), .S(n12609), .Y(n9789) );
  MUX2X1 U9410 ( .B(n9793), .A(n9794), .S(n12614), .Y(n9792) );
  MUX2X1 U9411 ( .B(n9796), .A(n9797), .S(mem_access_addr[3]), .Y(n9795) );
  MUX2X1 U9412 ( .B(n9799), .A(n9800), .S(n12592), .Y(n9798) );
  MUX2X1 U9413 ( .B(n9802), .A(n9803), .S(n12618), .Y(n9801) );
  MUX2X1 U9414 ( .B(n9805), .A(n9806), .S(n12596), .Y(n9804) );
  MUX2X1 U9415 ( .B(n9808), .A(n9809), .S(n12619), .Y(n9807) );
  MUX2X1 U9416 ( .B(n9811), .A(n9812), .S(n12572), .Y(n9810) );
  MUX2X1 U9417 ( .B(n9814), .A(n9815), .S(n12590), .Y(n9813) );
  MUX2X1 U9418 ( .B(n9817), .A(n9818), .S(n12619), .Y(n9816) );
  MUX2X1 U9419 ( .B(n9820), .A(n9821), .S(n12610), .Y(n9819) );
  MUX2X1 U9420 ( .B(n9823), .A(n9824), .S(n12617), .Y(n9822) );
  MUX2X1 U9421 ( .B(n9826), .A(n9827), .S(mem_access_addr[3]), .Y(n9825) );
  MUX2X1 U9422 ( .B(n9829), .A(n9830), .S(n12563), .Y(n9828) );
  MUX2X1 U9423 ( .B(n9832), .A(n9833), .S(n12616), .Y(n9831) );
  MUX2X1 U9424 ( .B(n9835), .A(n9836), .S(mem_access_addr[1]), .Y(n9834) );
  MUX2X1 U9425 ( .B(n9838), .A(n9839), .S(n12591), .Y(n9837) );
  MUX2X1 U9426 ( .B(n9841), .A(n9842), .S(n12596), .Y(n9840) );
  MUX2X1 U9427 ( .B(n9844), .A(n9845), .S(mem_access_addr[3]), .Y(n9843) );
  MUX2X1 U9428 ( .B(n9847), .A(n9848), .S(n12604), .Y(n9846) );
  MUX2X1 U9429 ( .B(n9850), .A(n9851), .S(n12599), .Y(n9849) );
  MUX2X1 U9430 ( .B(n9853), .A(n9854), .S(n12610), .Y(n9852) );
  MUX2X1 U9431 ( .B(n9856), .A(n9857), .S(n12593), .Y(n9855) );
  MUX2X1 U9432 ( .B(n9859), .A(n9860), .S(n12570), .Y(n9858) );
  MUX2X1 U9433 ( .B(n9862), .A(n9863), .S(n12608), .Y(n9861) );
  MUX2X1 U9434 ( .B(n9865), .A(n9866), .S(n12610), .Y(n9864) );
  MUX2X1 U9435 ( .B(n9868), .A(n9869), .S(n12603), .Y(n9867) );
  MUX2X1 U9436 ( .B(n9871), .A(n9872), .S(n12605), .Y(n9870) );
  MUX2X1 U9437 ( .B(n9874), .A(n9875), .S(mem_access_addr[3]), .Y(n9873) );
  MUX2X1 U9438 ( .B(n9877), .A(n9878), .S(n12618), .Y(n9876) );
  MUX2X1 U9439 ( .B(n9880), .A(n9881), .S(n12591), .Y(n9879) );
  MUX2X1 U9440 ( .B(n9883), .A(n9884), .S(n12608), .Y(n9882) );
  MUX2X1 U9441 ( .B(n9886), .A(n9887), .S(n12620), .Y(n9885) );
  MUX2X1 U9442 ( .B(n9889), .A(n9890), .S(n12574), .Y(n9888) );
  MUX2X1 U9443 ( .B(n9892), .A(n9893), .S(n12563), .Y(n9891) );
  MUX2X1 U9444 ( .B(n9895), .A(n9896), .S(n12593), .Y(n9894) );
  MUX2X1 U9445 ( .B(n9898), .A(n9899), .S(n12591), .Y(n9897) );
  MUX2X1 U9446 ( .B(n9901), .A(n9902), .S(n12593), .Y(n9900) );
  MUX2X1 U9447 ( .B(n9904), .A(n9905), .S(n12592), .Y(n9903) );
  MUX2X1 U9448 ( .B(n9907), .A(n9908), .S(n12570), .Y(n9906) );
  MUX2X1 U9449 ( .B(n9910), .A(n9911), .S(n12619), .Y(n9909) );
  MUX2X1 U9450 ( .B(n9913), .A(n9914), .S(n12614), .Y(n9912) );
  MUX2X1 U9451 ( .B(n9916), .A(n9917), .S(n12600), .Y(n9915) );
  MUX2X1 U9452 ( .B(n9919), .A(n9920), .S(n12603), .Y(n9918) );
  MUX2X1 U9453 ( .B(n9922), .A(n9923), .S(mem_access_addr[3]), .Y(n9921) );
  MUX2X1 U9454 ( .B(n9925), .A(n9926), .S(n12592), .Y(n9924) );
  MUX2X1 U9455 ( .B(n9928), .A(n9929), .S(n12612), .Y(n9927) );
  MUX2X1 U9456 ( .B(n9931), .A(n9932), .S(n12604), .Y(n9930) );
  MUX2X1 U9457 ( .B(n9934), .A(n9935), .S(n12604), .Y(n9933) );
  MUX2X1 U9458 ( .B(n9937), .A(n9938), .S(n12570), .Y(n9936) );
  MUX2X1 U9459 ( .B(n9940), .A(n9941), .S(n12618), .Y(n9939) );
  MUX2X1 U9460 ( .B(n9943), .A(n9944), .S(mem_access_addr[1]), .Y(n9942) );
  MUX2X1 U9461 ( .B(n9946), .A(n9947), .S(n12596), .Y(n9945) );
  MUX2X1 U9462 ( .B(n9949), .A(n9950), .S(n12592), .Y(n9948) );
  MUX2X1 U9463 ( .B(n9952), .A(n9953), .S(n12574), .Y(n9951) );
  MUX2X1 U9464 ( .B(n9955), .A(n9956), .S(n12562), .Y(n9954) );
  MUX2X1 U9465 ( .B(n9958), .A(n9959), .S(n12619), .Y(n9957) );
  MUX2X1 U9466 ( .B(n9961), .A(n9962), .S(mem_access_addr[1]), .Y(n9960) );
  MUX2X1 U9467 ( .B(n9964), .A(n9965), .S(n12596), .Y(n9963) );
  MUX2X1 U9468 ( .B(n9967), .A(n9968), .S(mem_access_addr[1]), .Y(n9966) );
  MUX2X1 U9469 ( .B(n9970), .A(n9971), .S(mem_access_addr[3]), .Y(n9969) );
  MUX2X1 U9470 ( .B(n9973), .A(n9974), .S(mem_access_addr[1]), .Y(n9972) );
  MUX2X1 U9471 ( .B(n9976), .A(n9977), .S(mem_access_addr[1]), .Y(n9975) );
  MUX2X1 U9472 ( .B(n9979), .A(n9980), .S(mem_access_addr[1]), .Y(n9978) );
  MUX2X1 U9473 ( .B(n9982), .A(n9983), .S(mem_access_addr[1]), .Y(n9981) );
  MUX2X1 U9474 ( .B(n9985), .A(n9986), .S(mem_access_addr[3]), .Y(n9984) );
  MUX2X1 U9475 ( .B(n9988), .A(n9989), .S(n12600), .Y(n9987) );
  MUX2X1 U9476 ( .B(n9991), .A(n9992), .S(n12610), .Y(n9990) );
  MUX2X1 U9477 ( .B(n9994), .A(n9995), .S(n12616), .Y(n9993) );
  MUX2X1 U9478 ( .B(n9997), .A(n9998), .S(n12590), .Y(n9996) );
  MUX2X1 U9479 ( .B(n10000), .A(n10001), .S(n12574), .Y(n9999) );
  MUX2X1 U9480 ( .B(n10003), .A(n10004), .S(n12596), .Y(n10002) );
  MUX2X1 U9481 ( .B(n10006), .A(n10007), .S(n12614), .Y(n10005) );
  MUX2X1 U9482 ( .B(n10009), .A(n10010), .S(n12595), .Y(n10008) );
  MUX2X1 U9483 ( .B(n10012), .A(n10013), .S(n12619), .Y(n10011) );
  MUX2X1 U9484 ( .B(n10015), .A(n10016), .S(mem_access_addr[3]), .Y(n10014) );
  MUX2X1 U9485 ( .B(n10018), .A(n10019), .S(n12563), .Y(n10017) );
  MUX2X1 U9486 ( .B(n10020), .A(n10021), .S(mem_access_addr[7]), .Y(
        mem_read_data[5]) );
  MUX2X1 U9487 ( .B(n10023), .A(n10024), .S(n12591), .Y(n10022) );
  MUX2X1 U9488 ( .B(n10026), .A(n10027), .S(n12620), .Y(n10025) );
  MUX2X1 U9489 ( .B(n10029), .A(n10030), .S(n12592), .Y(n10028) );
  MUX2X1 U9490 ( .B(n10032), .A(n10033), .S(n12605), .Y(n10031) );
  MUX2X1 U9491 ( .B(n10035), .A(n10036), .S(n12574), .Y(n10034) );
  MUX2X1 U9492 ( .B(n10038), .A(n10039), .S(n12604), .Y(n10037) );
  MUX2X1 U9493 ( .B(n10041), .A(n10042), .S(n12603), .Y(n10040) );
  MUX2X1 U9494 ( .B(n10044), .A(n10045), .S(n12611), .Y(n10043) );
  MUX2X1 U9495 ( .B(n10047), .A(n10048), .S(n12610), .Y(n10046) );
  MUX2X1 U9496 ( .B(n10050), .A(n10051), .S(mem_access_addr[3]), .Y(n10049) );
  MUX2X1 U9497 ( .B(n10053), .A(n10054), .S(n12615), .Y(n10052) );
  MUX2X1 U9498 ( .B(n10056), .A(n10057), .S(n12603), .Y(n10055) );
  MUX2X1 U9499 ( .B(n10059), .A(n10060), .S(n12593), .Y(n10058) );
  MUX2X1 U9500 ( .B(n10062), .A(n10063), .S(n12591), .Y(n10061) );
  MUX2X1 U9501 ( .B(n10065), .A(n10066), .S(n12574), .Y(n10064) );
  MUX2X1 U9502 ( .B(n10068), .A(n10069), .S(n12617), .Y(n10067) );
  MUX2X1 U9503 ( .B(n10071), .A(n10072), .S(n12618), .Y(n10070) );
  MUX2X1 U9504 ( .B(n10074), .A(n10075), .S(n12618), .Y(n10073) );
  MUX2X1 U9505 ( .B(n10077), .A(n10078), .S(n12590), .Y(n10076) );
  MUX2X1 U9506 ( .B(n10080), .A(n10081), .S(mem_access_addr[3]), .Y(n10079) );
  MUX2X1 U9507 ( .B(n10083), .A(n10084), .S(n12562), .Y(n10082) );
  MUX2X1 U9508 ( .B(n10086), .A(n10087), .S(n12620), .Y(n10085) );
  MUX2X1 U9509 ( .B(n10089), .A(n10090), .S(n12615), .Y(n10088) );
  MUX2X1 U9510 ( .B(n10092), .A(n10093), .S(n12601), .Y(n10091) );
  MUX2X1 U9511 ( .B(n10095), .A(n10096), .S(n12600), .Y(n10094) );
  MUX2X1 U9512 ( .B(n10098), .A(n10099), .S(n12572), .Y(n10097) );
  MUX2X1 U9513 ( .B(n10101), .A(n10102), .S(n12620), .Y(n10100) );
  MUX2X1 U9514 ( .B(n10104), .A(n10105), .S(n12619), .Y(n10103) );
  MUX2X1 U9515 ( .B(n10107), .A(n10108), .S(n12593), .Y(n10106) );
  MUX2X1 U9516 ( .B(n10110), .A(n10111), .S(n12601), .Y(n10109) );
  MUX2X1 U9517 ( .B(n10113), .A(n10114), .S(n12572), .Y(n10112) );
  MUX2X1 U9518 ( .B(n10116), .A(n10117), .S(n12596), .Y(n10115) );
  MUX2X1 U9519 ( .B(n10119), .A(n10120), .S(n12599), .Y(n10118) );
  MUX2X1 U9520 ( .B(n10122), .A(n10123), .S(n12602), .Y(n10121) );
  MUX2X1 U9521 ( .B(n10125), .A(n10126), .S(n12596), .Y(n10124) );
  MUX2X1 U9522 ( .B(n10128), .A(n10129), .S(n12568), .Y(n10127) );
  MUX2X1 U9523 ( .B(n10131), .A(n10132), .S(n12598), .Y(n10130) );
  MUX2X1 U9524 ( .B(n10134), .A(n10135), .S(n12613), .Y(n10133) );
  MUX2X1 U9525 ( .B(n10137), .A(n10138), .S(n12609), .Y(n10136) );
  MUX2X1 U9526 ( .B(n10140), .A(n10141), .S(n12602), .Y(n10139) );
  MUX2X1 U9527 ( .B(n10143), .A(n10144), .S(n12569), .Y(n10142) );
  MUX2X1 U9528 ( .B(n10146), .A(n10147), .S(n12562), .Y(n10145) );
  MUX2X1 U9529 ( .B(n10149), .A(n10150), .S(n12613), .Y(n10148) );
  MUX2X1 U9530 ( .B(n10152), .A(n10153), .S(n12620), .Y(n10151) );
  MUX2X1 U9531 ( .B(n10155), .A(n10156), .S(n12616), .Y(n10154) );
  MUX2X1 U9532 ( .B(n10158), .A(n10159), .S(n12603), .Y(n10157) );
  MUX2X1 U9533 ( .B(n10161), .A(n10162), .S(n12568), .Y(n10160) );
  MUX2X1 U9534 ( .B(n10164), .A(n10165), .S(n12608), .Y(n10163) );
  MUX2X1 U9535 ( .B(n10167), .A(n10168), .S(n12590), .Y(n10166) );
  MUX2X1 U9536 ( .B(n10170), .A(n10171), .S(n12597), .Y(n10169) );
  MUX2X1 U9537 ( .B(n10173), .A(n10174), .S(n12602), .Y(n10172) );
  MUX2X1 U9538 ( .B(n10176), .A(n10177), .S(n12572), .Y(n10175) );
  MUX2X1 U9539 ( .B(n10179), .A(n10180), .S(n12591), .Y(n10178) );
  MUX2X1 U9540 ( .B(n10182), .A(n10183), .S(n12597), .Y(n10181) );
  MUX2X1 U9541 ( .B(n10185), .A(n10186), .S(n12595), .Y(n10184) );
  MUX2X1 U9542 ( .B(n10188), .A(n10189), .S(n12618), .Y(n10187) );
  MUX2X1 U9543 ( .B(n10191), .A(n10192), .S(n12568), .Y(n10190) );
  MUX2X1 U9544 ( .B(n10194), .A(n10195), .S(n12604), .Y(n10193) );
  MUX2X1 U9545 ( .B(n10197), .A(n10198), .S(n12600), .Y(n10196) );
  MUX2X1 U9546 ( .B(n10200), .A(n10201), .S(n12605), .Y(n10199) );
  MUX2X1 U9547 ( .B(n10203), .A(n10204), .S(n12613), .Y(n10202) );
  MUX2X1 U9548 ( .B(n10206), .A(n10207), .S(n12572), .Y(n10205) );
  MUX2X1 U9549 ( .B(n10209), .A(n10210), .S(n12563), .Y(n10208) );
  MUX2X1 U9550 ( .B(n10212), .A(n10213), .S(n12596), .Y(n10211) );
  MUX2X1 U9551 ( .B(n10215), .A(n10216), .S(mem_access_addr[1]), .Y(n10214) );
  MUX2X1 U9552 ( .B(n10218), .A(n10219), .S(n12607), .Y(n10217) );
  MUX2X1 U9553 ( .B(n10221), .A(n10222), .S(n12601), .Y(n10220) );
  MUX2X1 U9554 ( .B(n10224), .A(n10225), .S(n12568), .Y(n10223) );
  MUX2X1 U9555 ( .B(n10227), .A(n10228), .S(n12606), .Y(n10226) );
  MUX2X1 U9556 ( .B(n10230), .A(n10231), .S(mem_access_addr[1]), .Y(n10229) );
  MUX2X1 U9557 ( .B(n10233), .A(n10234), .S(n12608), .Y(n10232) );
  MUX2X1 U9558 ( .B(n10236), .A(n10237), .S(n12604), .Y(n10235) );
  MUX2X1 U9559 ( .B(n10239), .A(n10240), .S(n12574), .Y(n10238) );
  MUX2X1 U9560 ( .B(n10242), .A(n10243), .S(n12608), .Y(n10241) );
  MUX2X1 U9561 ( .B(n10245), .A(n10246), .S(n12593), .Y(n10244) );
  MUX2X1 U9562 ( .B(n10248), .A(n10249), .S(n12598), .Y(n10247) );
  MUX2X1 U9563 ( .B(n10251), .A(n10252), .S(n12595), .Y(n10250) );
  MUX2X1 U9564 ( .B(n10254), .A(n10255), .S(n12570), .Y(n10253) );
  MUX2X1 U9565 ( .B(n10257), .A(n10258), .S(n12614), .Y(n10256) );
  MUX2X1 U9566 ( .B(n10260), .A(n10261), .S(n12592), .Y(n10259) );
  MUX2X1 U9567 ( .B(n10263), .A(n10264), .S(n12609), .Y(n10262) );
  MUX2X1 U9568 ( .B(n10266), .A(n10267), .S(n12611), .Y(n10265) );
  MUX2X1 U9569 ( .B(n10269), .A(n10270), .S(n12570), .Y(n10268) );
  MUX2X1 U9570 ( .B(n10272), .A(n10273), .S(n12562), .Y(n10271) );
  MUX2X1 U9571 ( .B(n10274), .A(n10275), .S(mem_access_addr[7]), .Y(
        mem_read_data[6]) );
  MUX2X1 U9572 ( .B(n10277), .A(n10278), .S(n12618), .Y(n10276) );
  MUX2X1 U9573 ( .B(n10280), .A(n10281), .S(n12590), .Y(n10279) );
  MUX2X1 U9574 ( .B(n10283), .A(n10284), .S(n12600), .Y(n10282) );
  MUX2X1 U9575 ( .B(n10286), .A(n10287), .S(n12602), .Y(n10285) );
  MUX2X1 U9576 ( .B(n10289), .A(n10290), .S(n12574), .Y(n10288) );
  MUX2X1 U9577 ( .B(n10292), .A(n10293), .S(n12609), .Y(n10291) );
  MUX2X1 U9578 ( .B(n10295), .A(n10296), .S(n12602), .Y(n10294) );
  MUX2X1 U9579 ( .B(n10298), .A(n10299), .S(n12617), .Y(n10297) );
  MUX2X1 U9580 ( .B(n10301), .A(n10302), .S(n12593), .Y(n10300) );
  MUX2X1 U9581 ( .B(n10304), .A(n10305), .S(mem_access_addr[3]), .Y(n10303) );
  MUX2X1 U9582 ( .B(n10307), .A(n10308), .S(n12596), .Y(n10306) );
  MUX2X1 U9583 ( .B(n10310), .A(n10311), .S(n12590), .Y(n10309) );
  MUX2X1 U9584 ( .B(n10313), .A(n10314), .S(n12594), .Y(n10312) );
  MUX2X1 U9585 ( .B(n10316), .A(n10317), .S(n12611), .Y(n10315) );
  MUX2X1 U9586 ( .B(n10319), .A(n10320), .S(n12570), .Y(n10318) );
  MUX2X1 U9587 ( .B(n10322), .A(n10323), .S(n12615), .Y(n10321) );
  MUX2X1 U9588 ( .B(n10325), .A(n10326), .S(n12615), .Y(n10324) );
  MUX2X1 U9589 ( .B(n10328), .A(n10329), .S(n12599), .Y(n10327) );
  MUX2X1 U9590 ( .B(n10331), .A(n10332), .S(n12615), .Y(n10330) );
  MUX2X1 U9591 ( .B(n10334), .A(n10335), .S(mem_access_addr[3]), .Y(n10333) );
  MUX2X1 U9592 ( .B(n10337), .A(n10338), .S(n12563), .Y(n10336) );
  MUX2X1 U9593 ( .B(n10340), .A(n10341), .S(n12595), .Y(n10339) );
  MUX2X1 U9594 ( .B(n10343), .A(n10344), .S(n12598), .Y(n10342) );
  MUX2X1 U9595 ( .B(n10346), .A(n10347), .S(n12609), .Y(n10345) );
  MUX2X1 U9596 ( .B(n10349), .A(n10350), .S(n12594), .Y(n10348) );
  MUX2X1 U9597 ( .B(n10352), .A(n10353), .S(mem_access_addr[3]), .Y(n10351) );
  MUX2X1 U9598 ( .B(n10355), .A(n10356), .S(n12617), .Y(n10354) );
  MUX2X1 U9599 ( .B(n10358), .A(n10359), .S(n12612), .Y(n10357) );
  MUX2X1 U9600 ( .B(n10361), .A(n10362), .S(n12612), .Y(n10360) );
  MUX2X1 U9601 ( .B(n10364), .A(n10365), .S(n12596), .Y(n10363) );
  MUX2X1 U9602 ( .B(n10367), .A(n10368), .S(mem_access_addr[3]), .Y(n10366) );
  MUX2X1 U9603 ( .B(n10370), .A(n10371), .S(n12591), .Y(n10369) );
  MUX2X1 U9604 ( .B(n10373), .A(n10374), .S(n12618), .Y(n10372) );
  MUX2X1 U9605 ( .B(n10376), .A(n10377), .S(n12605), .Y(n10375) );
  MUX2X1 U9606 ( .B(n10379), .A(n10380), .S(n12600), .Y(n10378) );
  MUX2X1 U9607 ( .B(n10382), .A(n10383), .S(mem_access_addr[3]), .Y(n10381) );
  MUX2X1 U9608 ( .B(n10385), .A(n10386), .S(mem_access_addr[1]), .Y(n10384) );
  MUX2X1 U9609 ( .B(n10388), .A(n10389), .S(n12612), .Y(n10387) );
  MUX2X1 U9610 ( .B(n10391), .A(n10392), .S(n12611), .Y(n10390) );
  MUX2X1 U9611 ( .B(n10394), .A(n10395), .S(n12613), .Y(n10393) );
  MUX2X1 U9612 ( .B(n10397), .A(n10398), .S(mem_access_addr[3]), .Y(n10396) );
  MUX2X1 U9613 ( .B(n10400), .A(n10401), .S(n12562), .Y(n10399) );
  MUX2X1 U9614 ( .B(n10403), .A(n10404), .S(n12606), .Y(n10402) );
  MUX2X1 U9615 ( .B(n10406), .A(n10407), .S(n12594), .Y(n10405) );
  MUX2X1 U9616 ( .B(n10409), .A(n10410), .S(n12595), .Y(n10408) );
  MUX2X1 U9617 ( .B(n10412), .A(n10413), .S(n12610), .Y(n10411) );
  MUX2X1 U9618 ( .B(n10415), .A(n10416), .S(n12571), .Y(n10414) );
  MUX2X1 U9619 ( .B(n10418), .A(n10419), .S(n12606), .Y(n10417) );
  MUX2X1 U9620 ( .B(n10421), .A(n10422), .S(n12591), .Y(n10420) );
  MUX2X1 U9621 ( .B(n10424), .A(n10425), .S(n12605), .Y(n10423) );
  MUX2X1 U9622 ( .B(n10427), .A(n10428), .S(n12614), .Y(n10426) );
  MUX2X1 U9623 ( .B(n10430), .A(n10431), .S(mem_access_addr[3]), .Y(n10429) );
  MUX2X1 U9624 ( .B(n10433), .A(n10434), .S(n12602), .Y(n10432) );
  MUX2X1 U9625 ( .B(n10436), .A(n10437), .S(n12590), .Y(n10435) );
  MUX2X1 U9626 ( .B(n10439), .A(n10440), .S(n12593), .Y(n10438) );
  MUX2X1 U9627 ( .B(n10442), .A(n10443), .S(n12602), .Y(n10441) );
  MUX2X1 U9628 ( .B(n10445), .A(n10446), .S(n12574), .Y(n10444) );
  MUX2X1 U9629 ( .B(n10448), .A(n10449), .S(n12593), .Y(n10447) );
  MUX2X1 U9630 ( .B(n10451), .A(n10452), .S(n12590), .Y(n10450) );
  MUX2X1 U9631 ( .B(n10454), .A(n10455), .S(n12603), .Y(n10453) );
  MUX2X1 U9632 ( .B(n10457), .A(n10458), .S(n12595), .Y(n10456) );
  MUX2X1 U9633 ( .B(n10460), .A(n10461), .S(n12574), .Y(n10459) );
  MUX2X1 U9634 ( .B(n10463), .A(n10464), .S(n12563), .Y(n10462) );
  MUX2X1 U9635 ( .B(n10466), .A(n10467), .S(n12593), .Y(n10465) );
  MUX2X1 U9636 ( .B(n10469), .A(n10470), .S(mem_access_addr[1]), .Y(n10468) );
  MUX2X1 U9637 ( .B(n10472), .A(n10473), .S(n12596), .Y(n10471) );
  MUX2X1 U9638 ( .B(n10475), .A(n10476), .S(mem_access_addr[1]), .Y(n10474) );
  MUX2X1 U9639 ( .B(n10478), .A(n10479), .S(mem_access_addr[3]), .Y(n10477) );
  MUX2X1 U9640 ( .B(n10481), .A(n10482), .S(mem_access_addr[1]), .Y(n10480) );
  MUX2X1 U9641 ( .B(n10484), .A(n10485), .S(mem_access_addr[1]), .Y(n10483) );
  MUX2X1 U9642 ( .B(n10487), .A(n10488), .S(mem_access_addr[1]), .Y(n10486) );
  MUX2X1 U9643 ( .B(n10490), .A(n10491), .S(mem_access_addr[1]), .Y(n10489) );
  MUX2X1 U9644 ( .B(n10493), .A(n10494), .S(n12574), .Y(n10492) );
  MUX2X1 U9645 ( .B(n10496), .A(n10497), .S(n12618), .Y(n10495) );
  MUX2X1 U9646 ( .B(n10499), .A(n10500), .S(mem_access_addr[1]), .Y(n10498) );
  MUX2X1 U9647 ( .B(n10502), .A(n10503), .S(n12603), .Y(n10501) );
  MUX2X1 U9648 ( .B(n10505), .A(n10506), .S(n12591), .Y(n10504) );
  MUX2X1 U9649 ( .B(n10508), .A(n10509), .S(n12572), .Y(n10507) );
  MUX2X1 U9650 ( .B(n10511), .A(n10512), .S(n12595), .Y(n10510) );
  MUX2X1 U9651 ( .B(n10514), .A(n10515), .S(n12607), .Y(n10513) );
  MUX2X1 U9652 ( .B(n10517), .A(n10518), .S(n12620), .Y(n10516) );
  MUX2X1 U9653 ( .B(n10520), .A(n10521), .S(n12592), .Y(n10519) );
  MUX2X1 U9654 ( .B(n10523), .A(n10524), .S(n12569), .Y(n10522) );
  MUX2X1 U9655 ( .B(n10526), .A(n10527), .S(n12563), .Y(n10525) );
  MUX2X1 U9656 ( .B(n10528), .A(n10529), .S(mem_access_addr[7]), .Y(
        mem_read_data[7]) );
  MUX2X1 U9657 ( .B(n10531), .A(n10532), .S(n12617), .Y(n10530) );
  MUX2X1 U9658 ( .B(n10534), .A(n10535), .S(n12613), .Y(n10533) );
  MUX2X1 U9659 ( .B(n10537), .A(n10538), .S(n12608), .Y(n10536) );
  MUX2X1 U9660 ( .B(n10540), .A(n10541), .S(n12597), .Y(n10539) );
  MUX2X1 U9661 ( .B(n10543), .A(n10544), .S(mem_access_addr[3]), .Y(n10542) );
  MUX2X1 U9662 ( .B(n10546), .A(n10547), .S(n12613), .Y(n10545) );
  MUX2X1 U9663 ( .B(n10549), .A(n10550), .S(n12609), .Y(n10548) );
  MUX2X1 U9664 ( .B(n10552), .A(n10553), .S(n12614), .Y(n10551) );
  MUX2X1 U9665 ( .B(n10555), .A(n10556), .S(mem_access_addr[1]), .Y(n10554) );
  MUX2X1 U9666 ( .B(n10558), .A(n10559), .S(n12571), .Y(n10557) );
  MUX2X1 U9667 ( .B(n10561), .A(n10562), .S(n12598), .Y(n10560) );
  MUX2X1 U9668 ( .B(n10564), .A(n10565), .S(n12609), .Y(n10563) );
  MUX2X1 U9669 ( .B(n10567), .A(n10568), .S(n12611), .Y(n10566) );
  MUX2X1 U9670 ( .B(n10570), .A(n10571), .S(n12594), .Y(n10569) );
  MUX2X1 U9671 ( .B(n10573), .A(n10574), .S(n12568), .Y(n10572) );
  MUX2X1 U9672 ( .B(n10576), .A(n10577), .S(n12597), .Y(n10575) );
  MUX2X1 U9673 ( .B(n10579), .A(n10580), .S(n12620), .Y(n10578) );
  MUX2X1 U9674 ( .B(n10582), .A(n10583), .S(n12610), .Y(n10581) );
  MUX2X1 U9675 ( .B(n10585), .A(n10586), .S(n12598), .Y(n10584) );
  MUX2X1 U9676 ( .B(n10588), .A(n10589), .S(n12574), .Y(n10587) );
  MUX2X1 U9677 ( .B(n10591), .A(n10592), .S(n12563), .Y(n10590) );
  MUX2X1 U9678 ( .B(n10594), .A(n10595), .S(n12618), .Y(n10593) );
  MUX2X1 U9679 ( .B(n10597), .A(n10598), .S(n12610), .Y(n10596) );
  MUX2X1 U9680 ( .B(n10600), .A(n10601), .S(n12608), .Y(n10599) );
  MUX2X1 U9681 ( .B(n10603), .A(n10604), .S(n12616), .Y(n10602) );
  MUX2X1 U9682 ( .B(n10606), .A(n10607), .S(mem_access_addr[3]), .Y(n10605) );
  MUX2X1 U9683 ( .B(n10609), .A(n10610), .S(n12620), .Y(n10608) );
  MUX2X1 U9684 ( .B(n10612), .A(n10613), .S(n12598), .Y(n10611) );
  MUX2X1 U9685 ( .B(n10615), .A(n10616), .S(n12620), .Y(n10614) );
  MUX2X1 U9686 ( .B(n10618), .A(n10619), .S(n12614), .Y(n10617) );
  MUX2X1 U9687 ( .B(n10621), .A(n10622), .S(n12574), .Y(n10620) );
  MUX2X1 U9688 ( .B(n10624), .A(n10625), .S(n12618), .Y(n10623) );
  MUX2X1 U9689 ( .B(n10627), .A(n10628), .S(n12619), .Y(n10626) );
  MUX2X1 U9690 ( .B(n10630), .A(n10631), .S(n12620), .Y(n10629) );
  MUX2X1 U9691 ( .B(n10633), .A(n10634), .S(n12618), .Y(n10632) );
  MUX2X1 U9692 ( .B(n10636), .A(n10637), .S(n12572), .Y(n10635) );
  MUX2X1 U9693 ( .B(n10639), .A(n10640), .S(n12619), .Y(n10638) );
  MUX2X1 U9694 ( .B(n10642), .A(n10643), .S(n12619), .Y(n10641) );
  MUX2X1 U9695 ( .B(n10645), .A(n10646), .S(n12590), .Y(n10644) );
  MUX2X1 U9696 ( .B(n10648), .A(n10649), .S(n12619), .Y(n10647) );
  MUX2X1 U9697 ( .B(n10651), .A(n10652), .S(n12570), .Y(n10650) );
  MUX2X1 U9698 ( .B(n10654), .A(n10655), .S(n12563), .Y(n10653) );
  MUX2X1 U9699 ( .B(n10657), .A(n10658), .S(n12608), .Y(n10656) );
  MUX2X1 U9700 ( .B(n10660), .A(n10661), .S(n12598), .Y(n10659) );
  MUX2X1 U9701 ( .B(n10663), .A(n10664), .S(n12594), .Y(n10662) );
  MUX2X1 U9702 ( .B(n10666), .A(n10667), .S(n12594), .Y(n10665) );
  MUX2X1 U9703 ( .B(n10669), .A(n10670), .S(n12568), .Y(n10668) );
  MUX2X1 U9704 ( .B(n10672), .A(n10673), .S(n12597), .Y(n10671) );
  MUX2X1 U9705 ( .B(n10675), .A(n10676), .S(n12594), .Y(n10674) );
  MUX2X1 U9706 ( .B(n10678), .A(n10679), .S(n12595), .Y(n10677) );
  MUX2X1 U9707 ( .B(n10681), .A(n10682), .S(n12605), .Y(n10680) );
  MUX2X1 U9708 ( .B(n10684), .A(n10685), .S(n12568), .Y(n10683) );
  MUX2X1 U9709 ( .B(n10687), .A(n10688), .S(n12608), .Y(n10686) );
  MUX2X1 U9710 ( .B(n10690), .A(n10691), .S(n12615), .Y(n10689) );
  MUX2X1 U9711 ( .B(n10693), .A(n10694), .S(n12610), .Y(n10692) );
  MUX2X1 U9712 ( .B(n10696), .A(n10697), .S(n12599), .Y(n10695) );
  MUX2X1 U9713 ( .B(n10699), .A(n10700), .S(n12568), .Y(n10698) );
  MUX2X1 U9714 ( .B(n10702), .A(n10703), .S(n12614), .Y(n10701) );
  MUX2X1 U9715 ( .B(n10705), .A(n10706), .S(n12607), .Y(n10704) );
  MUX2X1 U9716 ( .B(n10708), .A(n10709), .S(n12616), .Y(n10707) );
  MUX2X1 U9717 ( .B(n10711), .A(n10712), .S(n12618), .Y(n10710) );
  MUX2X1 U9718 ( .B(n10714), .A(n10715), .S(n12568), .Y(n10713) );
  MUX2X1 U9719 ( .B(n10717), .A(n10718), .S(n12562), .Y(n10716) );
  MUX2X1 U9720 ( .B(n10720), .A(n10721), .S(n12602), .Y(n10719) );
  MUX2X1 U9721 ( .B(n10723), .A(n10724), .S(n12596), .Y(n10722) );
  MUX2X1 U9722 ( .B(n10726), .A(n10727), .S(n12613), .Y(n10725) );
  MUX2X1 U9723 ( .B(n10729), .A(n10730), .S(n12616), .Y(n10728) );
  MUX2X1 U9724 ( .B(n10732), .A(n10733), .S(n12568), .Y(n10731) );
  MUX2X1 U9725 ( .B(n10735), .A(n10736), .S(n12611), .Y(n10734) );
  MUX2X1 U9726 ( .B(n10738), .A(n10739), .S(n12605), .Y(n10737) );
  MUX2X1 U9727 ( .B(n10741), .A(n10742), .S(n12593), .Y(n10740) );
  MUX2X1 U9728 ( .B(n10744), .A(n10745), .S(n12618), .Y(n10743) );
  MUX2X1 U9729 ( .B(n10747), .A(n10748), .S(n12568), .Y(n10746) );
  MUX2X1 U9730 ( .B(n10750), .A(n10751), .S(n12599), .Y(n10749) );
  MUX2X1 U9731 ( .B(n10753), .A(n10754), .S(n12614), .Y(n10752) );
  MUX2X1 U9732 ( .B(n10756), .A(n10757), .S(n12609), .Y(n10755) );
  MUX2X1 U9733 ( .B(n10759), .A(n10760), .S(n12592), .Y(n10758) );
  MUX2X1 U9734 ( .B(n10762), .A(n10763), .S(n12568), .Y(n10761) );
  MUX2X1 U9735 ( .B(n10765), .A(n10766), .S(n12600), .Y(n10764) );
  MUX2X1 U9736 ( .B(n10768), .A(n10769), .S(n12606), .Y(n10767) );
  MUX2X1 U9737 ( .B(n10771), .A(n10772), .S(n12611), .Y(n10770) );
  MUX2X1 U9738 ( .B(n10774), .A(n10775), .S(n12609), .Y(n10773) );
  MUX2X1 U9739 ( .B(n10777), .A(n10778), .S(n12568), .Y(n10776) );
  MUX2X1 U9740 ( .B(n10780), .A(n10781), .S(n12562), .Y(n10779) );
  MUX2X1 U9741 ( .B(n10782), .A(n10783), .S(mem_access_addr[7]), .Y(
        mem_read_data[8]) );
  MUX2X1 U9742 ( .B(n10785), .A(n10786), .S(n12614), .Y(n10784) );
  MUX2X1 U9743 ( .B(n10788), .A(n10789), .S(n12612), .Y(n10787) );
  MUX2X1 U9744 ( .B(n10791), .A(n10792), .S(n12608), .Y(n10790) );
  MUX2X1 U9745 ( .B(n10794), .A(n10795), .S(n12592), .Y(n10793) );
  MUX2X1 U9746 ( .B(n10797), .A(n10798), .S(n12568), .Y(n10796) );
  MUX2X1 U9747 ( .B(n10800), .A(n10801), .S(n12619), .Y(n10799) );
  MUX2X1 U9748 ( .B(n10803), .A(n10804), .S(n12610), .Y(n10802) );
  MUX2X1 U9749 ( .B(n10806), .A(n10807), .S(n12613), .Y(n10805) );
  MUX2X1 U9750 ( .B(n10809), .A(n10810), .S(n12597), .Y(n10808) );
  MUX2X1 U9751 ( .B(n10812), .A(n10813), .S(n12568), .Y(n10811) );
  MUX2X1 U9752 ( .B(n10815), .A(n10816), .S(n12615), .Y(n10814) );
  MUX2X1 U9753 ( .B(n10818), .A(n10819), .S(n12617), .Y(n10817) );
  MUX2X1 U9754 ( .B(n10821), .A(n10822), .S(n12605), .Y(n10820) );
  MUX2X1 U9755 ( .B(n10824), .A(n10825), .S(n12607), .Y(n10823) );
  MUX2X1 U9756 ( .B(n10827), .A(n10828), .S(n12568), .Y(n10826) );
  MUX2X1 U9757 ( .B(n10830), .A(n10831), .S(n12590), .Y(n10829) );
  MUX2X1 U9758 ( .B(n10833), .A(n10834), .S(n12604), .Y(n10832) );
  MUX2X1 U9759 ( .B(n10836), .A(n10837), .S(n12601), .Y(n10835) );
  MUX2X1 U9760 ( .B(n10839), .A(n10840), .S(n12596), .Y(n10838) );
  MUX2X1 U9761 ( .B(n10842), .A(n10843), .S(n12568), .Y(n10841) );
  MUX2X1 U9762 ( .B(n10845), .A(n10846), .S(n12562), .Y(n10844) );
  MUX2X1 U9763 ( .B(n10848), .A(n10849), .S(mem_access_addr[1]), .Y(n10847) );
  MUX2X1 U9764 ( .B(n10851), .A(n10852), .S(n12619), .Y(n10850) );
  MUX2X1 U9765 ( .B(n10854), .A(n10855), .S(n12594), .Y(n10853) );
  MUX2X1 U9766 ( .B(n10857), .A(n10858), .S(mem_access_addr[1]), .Y(n10856) );
  MUX2X1 U9767 ( .B(n10860), .A(n10861), .S(n12569), .Y(n10859) );
  MUX2X1 U9768 ( .B(n10863), .A(n10864), .S(n12620), .Y(n10862) );
  MUX2X1 U9769 ( .B(n10866), .A(n10867), .S(n12620), .Y(n10865) );
  MUX2X1 U9770 ( .B(n10869), .A(n10870), .S(mem_access_addr[1]), .Y(n10868) );
  MUX2X1 U9771 ( .B(n10872), .A(n10873), .S(n12618), .Y(n10871) );
  MUX2X1 U9772 ( .B(n10875), .A(n10876), .S(n12569), .Y(n10874) );
  MUX2X1 U9773 ( .B(n10878), .A(n10879), .S(n12610), .Y(n10877) );
  MUX2X1 U9774 ( .B(n10881), .A(n10882), .S(n12595), .Y(n10880) );
  MUX2X1 U9775 ( .B(n10884), .A(n10885), .S(n12596), .Y(n10883) );
  MUX2X1 U9776 ( .B(n10887), .A(n10888), .S(n12619), .Y(n10886) );
  MUX2X1 U9777 ( .B(n10890), .A(n10891), .S(n12569), .Y(n10889) );
  MUX2X1 U9778 ( .B(n10893), .A(n10894), .S(n12612), .Y(n10892) );
  MUX2X1 U9779 ( .B(n10896), .A(n10897), .S(n12590), .Y(n10895) );
  MUX2X1 U9780 ( .B(n10899), .A(n10900), .S(n12590), .Y(n10898) );
  MUX2X1 U9781 ( .B(n10902), .A(n10903), .S(n12618), .Y(n10901) );
  MUX2X1 U9782 ( .B(n10905), .A(n10906), .S(n12569), .Y(n10904) );
  MUX2X1 U9783 ( .B(n10908), .A(n10909), .S(n12563), .Y(n10907) );
  MUX2X1 U9784 ( .B(n10911), .A(n10912), .S(n12590), .Y(n10910) );
  MUX2X1 U9785 ( .B(n10914), .A(n10915), .S(n12593), .Y(n10913) );
  MUX2X1 U9786 ( .B(n10917), .A(n10918), .S(n12612), .Y(n10916) );
  MUX2X1 U9787 ( .B(n10920), .A(n10921), .S(n12617), .Y(n10919) );
  MUX2X1 U9788 ( .B(n10923), .A(n10924), .S(n12569), .Y(n10922) );
  MUX2X1 U9789 ( .B(n10926), .A(n10927), .S(n12619), .Y(n10925) );
  MUX2X1 U9790 ( .B(n10929), .A(n10930), .S(n12595), .Y(n10928) );
  MUX2X1 U9791 ( .B(n10932), .A(n10933), .S(n12592), .Y(n10931) );
  MUX2X1 U9792 ( .B(n10935), .A(n10936), .S(n12590), .Y(n10934) );
  MUX2X1 U9793 ( .B(n10938), .A(n10939), .S(n12569), .Y(n10937) );
  MUX2X1 U9794 ( .B(n10941), .A(n10942), .S(n12598), .Y(n10940) );
  MUX2X1 U9795 ( .B(n10944), .A(n10945), .S(n12593), .Y(n10943) );
  MUX2X1 U9796 ( .B(n10947), .A(n10948), .S(n12599), .Y(n10946) );
  MUX2X1 U9797 ( .B(n10950), .A(n10951), .S(n12596), .Y(n10949) );
  MUX2X1 U9798 ( .B(n10953), .A(n10954), .S(n12569), .Y(n10952) );
  MUX2X1 U9799 ( .B(n10956), .A(n10957), .S(n12595), .Y(n10955) );
  MUX2X1 U9800 ( .B(n10959), .A(n10960), .S(n12620), .Y(n10958) );
  MUX2X1 U9801 ( .B(n10962), .A(n10963), .S(n12601), .Y(n10961) );
  MUX2X1 U9802 ( .B(n10965), .A(n10966), .S(n12612), .Y(n10964) );
  MUX2X1 U9803 ( .B(n10968), .A(n10969), .S(n12569), .Y(n10967) );
  MUX2X1 U9804 ( .B(n10971), .A(n10972), .S(n12562), .Y(n10970) );
  MUX2X1 U9805 ( .B(n10974), .A(n10975), .S(n12616), .Y(n10973) );
  MUX2X1 U9806 ( .B(n10977), .A(n10978), .S(n12612), .Y(n10976) );
  MUX2X1 U9807 ( .B(n10980), .A(n10981), .S(n12603), .Y(n10979) );
  MUX2X1 U9808 ( .B(n10983), .A(n10984), .S(n12590), .Y(n10982) );
  MUX2X1 U9809 ( .B(n10986), .A(n10987), .S(n12569), .Y(n10985) );
  MUX2X1 U9810 ( .B(n10989), .A(n10990), .S(n12620), .Y(n10988) );
  MUX2X1 U9811 ( .B(n10992), .A(n10993), .S(n12603), .Y(n10991) );
  MUX2X1 U9812 ( .B(n10995), .A(n10996), .S(n12620), .Y(n10994) );
  MUX2X1 U9813 ( .B(n10998), .A(n10999), .S(n12594), .Y(n10997) );
  MUX2X1 U9814 ( .B(n11001), .A(n11002), .S(n12569), .Y(n11000) );
  MUX2X1 U9815 ( .B(n11004), .A(n11005), .S(n12599), .Y(n11003) );
  MUX2X1 U9816 ( .B(n11007), .A(n11008), .S(n12619), .Y(n11006) );
  MUX2X1 U9817 ( .B(n11010), .A(n11011), .S(n12600), .Y(n11009) );
  MUX2X1 U9818 ( .B(n11013), .A(n11014), .S(n12616), .Y(n11012) );
  MUX2X1 U9819 ( .B(n11016), .A(n11017), .S(n12569), .Y(n11015) );
  MUX2X1 U9820 ( .B(n11019), .A(n11020), .S(n12611), .Y(n11018) );
  MUX2X1 U9821 ( .B(n11022), .A(n11023), .S(n12592), .Y(n11021) );
  MUX2X1 U9822 ( .B(n11025), .A(n11026), .S(n12595), .Y(n11024) );
  MUX2X1 U9823 ( .B(n11028), .A(n11029), .S(n12615), .Y(n11027) );
  MUX2X1 U9824 ( .B(n11031), .A(n11032), .S(n12569), .Y(n11030) );
  MUX2X1 U9825 ( .B(n11034), .A(n11035), .S(n12563), .Y(n11033) );
  MUX2X1 U9826 ( .B(n11036), .A(n11037), .S(mem_access_addr[7]), .Y(
        mem_read_data[9]) );
  MUX2X1 U9827 ( .B(n11039), .A(n11040), .S(n12600), .Y(n11038) );
  MUX2X1 U9828 ( .B(n11042), .A(n11043), .S(n12592), .Y(n11041) );
  MUX2X1 U9829 ( .B(n11045), .A(n11046), .S(n12612), .Y(n11044) );
  MUX2X1 U9830 ( .B(n11048), .A(n11049), .S(n12605), .Y(n11047) );
  MUX2X1 U9831 ( .B(n11051), .A(n11052), .S(n12570), .Y(n11050) );
  MUX2X1 U9832 ( .B(n11054), .A(n11055), .S(n12594), .Y(n11053) );
  MUX2X1 U9833 ( .B(n11057), .A(n11058), .S(n12591), .Y(n11056) );
  MUX2X1 U9834 ( .B(n11060), .A(n11061), .S(n12607), .Y(n11059) );
  MUX2X1 U9835 ( .B(n11063), .A(n11064), .S(n12618), .Y(n11062) );
  MUX2X1 U9836 ( .B(n11066), .A(n11067), .S(n12570), .Y(n11065) );
  MUX2X1 U9837 ( .B(n11069), .A(n11070), .S(n12595), .Y(n11068) );
  MUX2X1 U9838 ( .B(n11072), .A(n11073), .S(n12596), .Y(n11071) );
  MUX2X1 U9839 ( .B(n11075), .A(n11076), .S(n12609), .Y(n11074) );
  MUX2X1 U9840 ( .B(n11078), .A(n11079), .S(n12608), .Y(n11077) );
  MUX2X1 U9841 ( .B(n11081), .A(n11082), .S(n12570), .Y(n11080) );
  MUX2X1 U9842 ( .B(n11084), .A(n11085), .S(n12595), .Y(n11083) );
  MUX2X1 U9843 ( .B(n11087), .A(n11088), .S(n12591), .Y(n11086) );
  MUX2X1 U9844 ( .B(n11090), .A(n11091), .S(n12594), .Y(n11089) );
  MUX2X1 U9845 ( .B(n11093), .A(n11094), .S(n12619), .Y(n11092) );
  MUX2X1 U9846 ( .B(n11096), .A(n11097), .S(n12570), .Y(n11095) );
  MUX2X1 U9847 ( .B(n11099), .A(n11100), .S(n12563), .Y(n11098) );
  MUX2X1 U9848 ( .B(n11102), .A(n11103), .S(n12603), .Y(n11101) );
  MUX2X1 U9849 ( .B(n11105), .A(n11106), .S(n12608), .Y(n11104) );
  MUX2X1 U9850 ( .B(n11108), .A(n11109), .S(n12613), .Y(n11107) );
  MUX2X1 U9851 ( .B(n11111), .A(n11112), .S(n12591), .Y(n11110) );
  MUX2X1 U9852 ( .B(n11114), .A(n11115), .S(n12570), .Y(n11113) );
  MUX2X1 U9853 ( .B(n11117), .A(n11118), .S(n12599), .Y(n11116) );
  MUX2X1 U9854 ( .B(n11120), .A(n11121), .S(n12606), .Y(n11119) );
  MUX2X1 U9855 ( .B(n11123), .A(n11124), .S(n12619), .Y(n11122) );
  MUX2X1 U9856 ( .B(n11126), .A(n11127), .S(n12602), .Y(n11125) );
  MUX2X1 U9857 ( .B(n11129), .A(n11130), .S(n12570), .Y(n11128) );
  MUX2X1 U9858 ( .B(n11132), .A(n11133), .S(n12596), .Y(n11131) );
  MUX2X1 U9859 ( .B(n11135), .A(n11136), .S(n12620), .Y(n11134) );
  MUX2X1 U9860 ( .B(n11138), .A(n11139), .S(n12607), .Y(n11137) );
  MUX2X1 U9861 ( .B(n11141), .A(n11142), .S(n12606), .Y(n11140) );
  MUX2X1 U9862 ( .B(n11144), .A(n11145), .S(n12570), .Y(n11143) );
  MUX2X1 U9863 ( .B(n11147), .A(n11148), .S(n12601), .Y(n11146) );
  MUX2X1 U9864 ( .B(n11150), .A(n11151), .S(n12607), .Y(n11149) );
  MUX2X1 U9865 ( .B(n11153), .A(n11154), .S(n12604), .Y(n11152) );
  MUX2X1 U9866 ( .B(n11156), .A(n11157), .S(n12591), .Y(n11155) );
  MUX2X1 U9867 ( .B(n11159), .A(n11160), .S(n12570), .Y(n11158) );
  MUX2X1 U9868 ( .B(n11162), .A(n11163), .S(n12563), .Y(n11161) );
  MUX2X1 U9869 ( .B(n11165), .A(n11166), .S(n12606), .Y(n11164) );
  MUX2X1 U9870 ( .B(n11168), .A(n11169), .S(n12611), .Y(n11167) );
  MUX2X1 U9871 ( .B(n11171), .A(n11172), .S(n12599), .Y(n11170) );
  MUX2X1 U9872 ( .B(n11174), .A(n11175), .S(n12616), .Y(n11173) );
  MUX2X1 U9873 ( .B(n11177), .A(n11178), .S(n12570), .Y(n11176) );
  MUX2X1 U9874 ( .B(n11180), .A(n11181), .S(n12618), .Y(n11179) );
  MUX2X1 U9875 ( .B(n11183), .A(n11184), .S(n12594), .Y(n11182) );
  MUX2X1 U9876 ( .B(n11186), .A(n11187), .S(n12616), .Y(n11185) );
  MUX2X1 U9877 ( .B(n11189), .A(n11190), .S(n12617), .Y(n11188) );
  MUX2X1 U9878 ( .B(n11192), .A(n11193), .S(n12570), .Y(n11191) );
  MUX2X1 U9879 ( .B(n11195), .A(n11196), .S(n12601), .Y(n11194) );
  MUX2X1 U9880 ( .B(n11198), .A(n11199), .S(n12608), .Y(n11197) );
  MUX2X1 U9881 ( .B(n11201), .A(n11202), .S(n12613), .Y(n11200) );
  MUX2X1 U9882 ( .B(n11204), .A(n11205), .S(n12615), .Y(n11203) );
  MUX2X1 U9883 ( .B(n11207), .A(n11208), .S(n12570), .Y(n11206) );
  MUX2X1 U9884 ( .B(n11210), .A(n11211), .S(n12597), .Y(n11209) );
  MUX2X1 U9885 ( .B(n11213), .A(n11214), .S(n12593), .Y(n11212) );
  MUX2X1 U9886 ( .B(n11216), .A(n11217), .S(n12610), .Y(n11215) );
  MUX2X1 U9887 ( .B(n11219), .A(n11220), .S(n12609), .Y(n11218) );
  MUX2X1 U9888 ( .B(n11222), .A(n11223), .S(n12570), .Y(n11221) );
  MUX2X1 U9889 ( .B(n11225), .A(n11226), .S(n12562), .Y(n11224) );
  MUX2X1 U9890 ( .B(n11228), .A(n11229), .S(n12614), .Y(n11227) );
  MUX2X1 U9891 ( .B(n11231), .A(n11232), .S(n12594), .Y(n11230) );
  MUX2X1 U9892 ( .B(n11234), .A(n11235), .S(n12592), .Y(n11233) );
  MUX2X1 U9893 ( .B(n11237), .A(n11238), .S(n12592), .Y(n11236) );
  MUX2X1 U9894 ( .B(n11240), .A(n11241), .S(n12569), .Y(n11239) );
  MUX2X1 U9895 ( .B(n11243), .A(n11244), .S(n12592), .Y(n11242) );
  MUX2X1 U9896 ( .B(n11246), .A(n11247), .S(n12616), .Y(n11245) );
  MUX2X1 U9897 ( .B(n11249), .A(n11250), .S(n12595), .Y(n11248) );
  MUX2X1 U9898 ( .B(n11252), .A(n11253), .S(n12593), .Y(n11251) );
  MUX2X1 U9899 ( .B(n11255), .A(n11256), .S(n12570), .Y(n11254) );
  MUX2X1 U9900 ( .B(n11258), .A(n11259), .S(n12590), .Y(n11257) );
  MUX2X1 U9901 ( .B(n11261), .A(n11262), .S(n12595), .Y(n11260) );
  MUX2X1 U9902 ( .B(n11264), .A(n11265), .S(n12600), .Y(n11263) );
  MUX2X1 U9903 ( .B(n11267), .A(n11268), .S(n12605), .Y(n11266) );
  MUX2X1 U9904 ( .B(n11270), .A(n11271), .S(n12574), .Y(n11269) );
  MUX2X1 U9905 ( .B(n11273), .A(n11274), .S(n12597), .Y(n11272) );
  MUX2X1 U9906 ( .B(n11276), .A(n11277), .S(n12597), .Y(n11275) );
  MUX2X1 U9907 ( .B(n11279), .A(n11280), .S(n12597), .Y(n11278) );
  MUX2X1 U9908 ( .B(n11282), .A(n11283), .S(n12597), .Y(n11281) );
  MUX2X1 U9909 ( .B(n11285), .A(n11286), .S(n12572), .Y(n11284) );
  MUX2X1 U9910 ( .B(n11288), .A(n11289), .S(n12562), .Y(n11287) );
  MUX2X1 U9911 ( .B(n11290), .A(n11291), .S(mem_access_addr[7]), .Y(
        mem_read_data[10]) );
  MUX2X1 U9912 ( .B(n11293), .A(n11294), .S(n12597), .Y(n11292) );
  MUX2X1 U9913 ( .B(n11296), .A(n11297), .S(n12597), .Y(n11295) );
  MUX2X1 U9914 ( .B(n11299), .A(n11300), .S(n12597), .Y(n11298) );
  MUX2X1 U9915 ( .B(n11302), .A(n11303), .S(n12597), .Y(n11301) );
  MUX2X1 U9916 ( .B(n11305), .A(n11306), .S(n12569), .Y(n11304) );
  MUX2X1 U9917 ( .B(n11308), .A(n11309), .S(n12597), .Y(n11307) );
  MUX2X1 U9918 ( .B(n11311), .A(n11312), .S(n12597), .Y(n11310) );
  MUX2X1 U9919 ( .B(n11314), .A(n11315), .S(n12597), .Y(n11313) );
  MUX2X1 U9920 ( .B(n11317), .A(n11318), .S(n12597), .Y(n11316) );
  MUX2X1 U9921 ( .B(n11320), .A(n11321), .S(n12571), .Y(n11319) );
  MUX2X1 U9922 ( .B(n11323), .A(n11324), .S(n12609), .Y(n11322) );
  MUX2X1 U9923 ( .B(n11326), .A(n11327), .S(n12594), .Y(n11325) );
  MUX2X1 U9924 ( .B(n11329), .A(n11330), .S(n12615), .Y(n11328) );
  MUX2X1 U9925 ( .B(n11332), .A(n11333), .S(n12599), .Y(n11331) );
  MUX2X1 U9926 ( .B(n11335), .A(n11336), .S(n12571), .Y(n11334) );
  MUX2X1 U9927 ( .B(n11338), .A(n11339), .S(n12612), .Y(n11337) );
  MUX2X1 U9928 ( .B(n11341), .A(n11342), .S(n12616), .Y(n11340) );
  MUX2X1 U9929 ( .B(n11344), .A(n11345), .S(n12600), .Y(n11343) );
  MUX2X1 U9930 ( .B(n11347), .A(n11348), .S(n12619), .Y(n11346) );
  MUX2X1 U9931 ( .B(n11350), .A(n11351), .S(n12571), .Y(n11349) );
  MUX2X1 U9932 ( .B(n11353), .A(n11354), .S(n12562), .Y(n11352) );
  MUX2X1 U9933 ( .B(n11356), .A(n11357), .S(n12596), .Y(n11355) );
  MUX2X1 U9934 ( .B(n11359), .A(n11360), .S(n12620), .Y(n11358) );
  MUX2X1 U9935 ( .B(n11362), .A(n11363), .S(n12593), .Y(n11361) );
  MUX2X1 U9936 ( .B(n11365), .A(n11366), .S(n12601), .Y(n11364) );
  MUX2X1 U9937 ( .B(n11368), .A(n11369), .S(n12569), .Y(n11367) );
  MUX2X1 U9938 ( .B(n11371), .A(n11372), .S(n12596), .Y(n11370) );
  MUX2X1 U9939 ( .B(n11374), .A(n11375), .S(n12610), .Y(n11373) );
  MUX2X1 U9940 ( .B(n11377), .A(n11378), .S(n12594), .Y(n11376) );
  MUX2X1 U9941 ( .B(n11380), .A(n11381), .S(n12594), .Y(n11379) );
  MUX2X1 U9942 ( .B(n11383), .A(n11384), .S(n12572), .Y(n11382) );
  MUX2X1 U9943 ( .B(n11386), .A(n11387), .S(n12593), .Y(n11385) );
  MUX2X1 U9944 ( .B(n11389), .A(n11390), .S(n12598), .Y(n11388) );
  MUX2X1 U9945 ( .B(n11392), .A(n11393), .S(n12591), .Y(n11391) );
  MUX2X1 U9946 ( .B(n11395), .A(n11396), .S(n12606), .Y(n11394) );
  MUX2X1 U9947 ( .B(n11398), .A(n11399), .S(n12570), .Y(n11397) );
  MUX2X1 U9948 ( .B(n11401), .A(n11402), .S(n12595), .Y(n11400) );
  MUX2X1 U9949 ( .B(n11404), .A(n11405), .S(n12611), .Y(n11403) );
  MUX2X1 U9950 ( .B(n11407), .A(n11408), .S(n12604), .Y(n11406) );
  MUX2X1 U9951 ( .B(n11410), .A(n11411), .S(n12602), .Y(n11409) );
  MUX2X1 U9952 ( .B(n11413), .A(n11414), .S(n12572), .Y(n11412) );
  MUX2X1 U9953 ( .B(n11416), .A(n11417), .S(n12562), .Y(n11415) );
  MUX2X1 U9954 ( .B(n11419), .A(n11420), .S(n12597), .Y(n11418) );
  MUX2X1 U9955 ( .B(n11422), .A(n11423), .S(n12592), .Y(n11421) );
  MUX2X1 U9956 ( .B(n11425), .A(n11426), .S(n12594), .Y(n11424) );
  MUX2X1 U9957 ( .B(n11428), .A(n11429), .S(n12606), .Y(n11427) );
  MUX2X1 U9958 ( .B(n11431), .A(n11432), .S(n12571), .Y(n11430) );
  MUX2X1 U9959 ( .B(n11434), .A(n11435), .S(n12615), .Y(n11433) );
  MUX2X1 U9960 ( .B(n11437), .A(n11438), .S(n12618), .Y(n11436) );
  MUX2X1 U9961 ( .B(n11440), .A(n11441), .S(n12611), .Y(n11439) );
  MUX2X1 U9962 ( .B(n11443), .A(n11444), .S(n12595), .Y(n11442) );
  MUX2X1 U9963 ( .B(n11446), .A(n11447), .S(n12574), .Y(n11445) );
  MUX2X1 U9964 ( .B(n11449), .A(n11450), .S(n12592), .Y(n11448) );
  MUX2X1 U9965 ( .B(n11452), .A(n11453), .S(n12593), .Y(n11451) );
  MUX2X1 U9966 ( .B(n11455), .A(n11456), .S(n12598), .Y(n11454) );
  MUX2X1 U9967 ( .B(n11458), .A(n11459), .S(n12590), .Y(n11457) );
  MUX2X1 U9968 ( .B(n11461), .A(n11462), .S(n12569), .Y(n11460) );
  MUX2X1 U9969 ( .B(n11464), .A(n11465), .S(n12599), .Y(n11463) );
  MUX2X1 U9970 ( .B(n11467), .A(n11468), .S(n12606), .Y(n11466) );
  MUX2X1 U9971 ( .B(n11470), .A(n11471), .S(n12602), .Y(n11469) );
  MUX2X1 U9972 ( .B(n11473), .A(n11474), .S(n12602), .Y(n11472) );
  MUX2X1 U9973 ( .B(n11476), .A(n11477), .S(n12571), .Y(n11475) );
  MUX2X1 U9974 ( .B(n11479), .A(n11480), .S(n12563), .Y(n11478) );
  MUX2X1 U9975 ( .B(n11482), .A(n11483), .S(n12590), .Y(n11481) );
  MUX2X1 U9976 ( .B(n11485), .A(n11486), .S(n12601), .Y(n11484) );
  MUX2X1 U9977 ( .B(n11488), .A(n11489), .S(n12611), .Y(n11487) );
  MUX2X1 U9978 ( .B(n11491), .A(n11492), .S(n12606), .Y(n11490) );
  MUX2X1 U9979 ( .B(n11494), .A(n11495), .S(n12574), .Y(n11493) );
  MUX2X1 U9980 ( .B(n11497), .A(n11498), .S(n12603), .Y(n11496) );
  MUX2X1 U9981 ( .B(n11500), .A(n11501), .S(n12617), .Y(n11499) );
  MUX2X1 U9982 ( .B(n11503), .A(n11504), .S(n12591), .Y(n11502) );
  MUX2X1 U9983 ( .B(n11506), .A(n11507), .S(n12596), .Y(n11505) );
  MUX2X1 U9984 ( .B(n11509), .A(n11510), .S(n12569), .Y(n11508) );
  MUX2X1 U9985 ( .B(n11512), .A(n11513), .S(n12598), .Y(n11511) );
  MUX2X1 U9986 ( .B(n11515), .A(n11516), .S(n12594), .Y(n11514) );
  MUX2X1 U9987 ( .B(n11518), .A(n11519), .S(n12615), .Y(n11517) );
  MUX2X1 U9988 ( .B(n11521), .A(n11522), .S(n12603), .Y(n11520) );
  MUX2X1 U9989 ( .B(n11524), .A(n11525), .S(n12572), .Y(n11523) );
  MUX2X1 U9990 ( .B(n11527), .A(n11528), .S(n12600), .Y(n11526) );
  MUX2X1 U9991 ( .B(n11530), .A(n11531), .S(n12596), .Y(n11529) );
  MUX2X1 U9992 ( .B(n11533), .A(n11534), .S(n12604), .Y(n11532) );
  MUX2X1 U9993 ( .B(n11536), .A(n11537), .S(n12590), .Y(n11535) );
  MUX2X1 U9994 ( .B(n11539), .A(n11540), .S(n12571), .Y(n11538) );
  MUX2X1 U9995 ( .B(n11542), .A(n11543), .S(n12563), .Y(n11541) );
  MUX2X1 U9996 ( .B(n11544), .A(n11545), .S(mem_access_addr[7]), .Y(
        mem_read_data[11]) );
  MUX2X1 U9997 ( .B(n11547), .A(n11548), .S(n12601), .Y(n11546) );
  MUX2X1 U9998 ( .B(n11550), .A(n11551), .S(n12620), .Y(n11549) );
  MUX2X1 U9999 ( .B(n11553), .A(n11554), .S(n12608), .Y(n11552) );
  MUX2X1 U10000 ( .B(n11556), .A(n11557), .S(n12593), .Y(n11555) );
  MUX2X1 U10001 ( .B(n11559), .A(n11560), .S(n12570), .Y(n11558) );
  MUX2X1 U10002 ( .B(n11562), .A(n11563), .S(n12613), .Y(n11561) );
  MUX2X1 U10003 ( .B(n11565), .A(n11566), .S(n12619), .Y(n11564) );
  MUX2X1 U10004 ( .B(n11568), .A(n11569), .S(n12616), .Y(n11567) );
  MUX2X1 U10005 ( .B(n11571), .A(n11572), .S(n12591), .Y(n11570) );
  MUX2X1 U10006 ( .B(n11574), .A(n11575), .S(n12572), .Y(n11573) );
  MUX2X1 U10007 ( .B(n11577), .A(n11578), .S(n12592), .Y(n11576) );
  MUX2X1 U10008 ( .B(n11580), .A(n11581), .S(n12607), .Y(n11579) );
  MUX2X1 U10009 ( .B(n11583), .A(n11584), .S(n12595), .Y(n11582) );
  MUX2X1 U10010 ( .B(n11586), .A(n11587), .S(n12599), .Y(n11585) );
  MUX2X1 U10011 ( .B(n11589), .A(n11590), .S(n12572), .Y(n11588) );
  MUX2X1 U10012 ( .B(n11592), .A(n11593), .S(n12620), .Y(n11591) );
  MUX2X1 U10013 ( .B(n11595), .A(n11596), .S(n12609), .Y(n11594) );
  MUX2X1 U10014 ( .B(n11598), .A(n11599), .S(n12600), .Y(n11597) );
  MUX2X1 U10015 ( .B(n11601), .A(n11602), .S(n12592), .Y(n11600) );
  MUX2X1 U10016 ( .B(n11604), .A(n11605), .S(n12574), .Y(n11603) );
  MUX2X1 U10017 ( .B(n11607), .A(n11608), .S(n12563), .Y(n11606) );
  MUX2X1 U10018 ( .B(n11610), .A(n11611), .S(n12598), .Y(n11609) );
  MUX2X1 U10019 ( .B(n11613), .A(n11614), .S(n12598), .Y(n11612) );
  MUX2X1 U10020 ( .B(n11616), .A(n11617), .S(n12598), .Y(n11615) );
  MUX2X1 U10021 ( .B(n11619), .A(n11620), .S(n12598), .Y(n11618) );
  MUX2X1 U10022 ( .B(n11622), .A(n11623), .S(n12569), .Y(n11621) );
  MUX2X1 U10023 ( .B(n11625), .A(n11626), .S(n12598), .Y(n11624) );
  MUX2X1 U10024 ( .B(n11628), .A(n11629), .S(n12598), .Y(n11627) );
  MUX2X1 U10025 ( .B(n11631), .A(n11632), .S(n12598), .Y(n11630) );
  MUX2X1 U10026 ( .B(n11634), .A(n11635), .S(n12598), .Y(n11633) );
  MUX2X1 U10027 ( .B(n11637), .A(n11638), .S(n12574), .Y(n11636) );
  MUX2X1 U10028 ( .B(n11640), .A(n11641), .S(n12598), .Y(n11639) );
  MUX2X1 U10029 ( .B(n11643), .A(n11644), .S(n12598), .Y(n11642) );
  MUX2X1 U10030 ( .B(n11646), .A(n11647), .S(n12598), .Y(n11645) );
  MUX2X1 U10031 ( .B(n11649), .A(n11650), .S(n12598), .Y(n11648) );
  MUX2X1 U10032 ( .B(n11652), .A(n11653), .S(n12569), .Y(n11651) );
  MUX2X1 U10033 ( .B(n11655), .A(n11656), .S(n12599), .Y(n11654) );
  MUX2X1 U10034 ( .B(n11658), .A(n11659), .S(n12599), .Y(n11657) );
  MUX2X1 U10035 ( .B(n11661), .A(n11662), .S(n12599), .Y(n11660) );
  MUX2X1 U10036 ( .B(n11664), .A(n11665), .S(n12599), .Y(n11663) );
  MUX2X1 U10037 ( .B(n11667), .A(n11668), .S(n12574), .Y(n11666) );
  MUX2X1 U10038 ( .B(n11670), .A(n11671), .S(n12562), .Y(n11669) );
  MUX2X1 U10039 ( .B(n11673), .A(n11674), .S(n12599), .Y(n11672) );
  MUX2X1 U10040 ( .B(n11676), .A(n11677), .S(n12599), .Y(n11675) );
  MUX2X1 U10041 ( .B(n11679), .A(n11680), .S(n12599), .Y(n11678) );
  MUX2X1 U10042 ( .B(n11682), .A(n11683), .S(n12599), .Y(n11681) );
  MUX2X1 U10043 ( .B(n11685), .A(n11686), .S(n12573), .Y(n11684) );
  MUX2X1 U10044 ( .B(n11688), .A(n11689), .S(n12599), .Y(n11687) );
  MUX2X1 U10045 ( .B(n11691), .A(n11692), .S(n12599), .Y(n11690) );
  MUX2X1 U10046 ( .B(n11694), .A(n11695), .S(n12599), .Y(n11693) );
  MUX2X1 U10047 ( .B(n11697), .A(n11698), .S(n12599), .Y(n11696) );
  MUX2X1 U10048 ( .B(n11700), .A(n11701), .S(n12572), .Y(n11699) );
  MUX2X1 U10049 ( .B(n11703), .A(n11704), .S(n12600), .Y(n11702) );
  MUX2X1 U10050 ( .B(n11706), .A(n11707), .S(n12600), .Y(n11705) );
  MUX2X1 U10051 ( .B(n11709), .A(n11710), .S(n12600), .Y(n11708) );
  MUX2X1 U10052 ( .B(n11712), .A(n11713), .S(n12600), .Y(n11711) );
  MUX2X1 U10053 ( .B(n11715), .A(n11716), .S(n12573), .Y(n11714) );
  MUX2X1 U10054 ( .B(n11718), .A(n11719), .S(n12600), .Y(n11717) );
  MUX2X1 U10055 ( .B(n11721), .A(n11722), .S(n12600), .Y(n11720) );
  MUX2X1 U10056 ( .B(n11724), .A(n11725), .S(n12600), .Y(n11723) );
  MUX2X1 U10057 ( .B(n11727), .A(n11728), .S(n12600), .Y(n11726) );
  MUX2X1 U10058 ( .B(n11730), .A(n11731), .S(n12569), .Y(n11729) );
  MUX2X1 U10059 ( .B(n11733), .A(n11734), .S(n12563), .Y(n11732) );
  MUX2X1 U10060 ( .B(n11736), .A(n11737), .S(n12600), .Y(n11735) );
  MUX2X1 U10061 ( .B(n11739), .A(n11740), .S(n12600), .Y(n11738) );
  MUX2X1 U10062 ( .B(n11742), .A(n11743), .S(n12600), .Y(n11741) );
  MUX2X1 U10063 ( .B(n11745), .A(n11746), .S(n12600), .Y(n11744) );
  MUX2X1 U10064 ( .B(n11748), .A(n11749), .S(n12570), .Y(n11747) );
  MUX2X1 U10065 ( .B(n11751), .A(n11752), .S(n12601), .Y(n11750) );
  MUX2X1 U10066 ( .B(n11754), .A(n11755), .S(n12601), .Y(n11753) );
  MUX2X1 U10067 ( .B(n11757), .A(n11758), .S(n12601), .Y(n11756) );
  MUX2X1 U10068 ( .B(n11760), .A(n11761), .S(n12601), .Y(n11759) );
  MUX2X1 U10069 ( .B(n11763), .A(n11764), .S(n12571), .Y(n11762) );
  MUX2X1 U10070 ( .B(n11766), .A(n11767), .S(n12601), .Y(n11765) );
  MUX2X1 U10071 ( .B(n11769), .A(n11770), .S(n12601), .Y(n11768) );
  MUX2X1 U10072 ( .B(n11772), .A(n11773), .S(n12601), .Y(n11771) );
  MUX2X1 U10073 ( .B(n11775), .A(n11776), .S(n12601), .Y(n11774) );
  MUX2X1 U10074 ( .B(n11778), .A(n11779), .S(n12572), .Y(n11777) );
  MUX2X1 U10075 ( .B(n11781), .A(n11782), .S(n12601), .Y(n11780) );
  MUX2X1 U10076 ( .B(n11784), .A(n11785), .S(n12601), .Y(n11783) );
  MUX2X1 U10077 ( .B(n11787), .A(n11788), .S(n12601), .Y(n11786) );
  MUX2X1 U10078 ( .B(n11790), .A(n11791), .S(n12601), .Y(n11789) );
  MUX2X1 U10079 ( .B(n11793), .A(n11794), .S(n12572), .Y(n11792) );
  MUX2X1 U10080 ( .B(n11796), .A(n11797), .S(n12562), .Y(n11795) );
  MUX2X1 U10081 ( .B(n11798), .A(n11799), .S(mem_access_addr[7]), .Y(
        mem_read_data[12]) );
  MUX2X1 U10082 ( .B(n11801), .A(n11802), .S(n12602), .Y(n11800) );
  MUX2X1 U10083 ( .B(n11804), .A(n11805), .S(n12602), .Y(n11803) );
  MUX2X1 U10084 ( .B(n11807), .A(n11808), .S(n12602), .Y(n11806) );
  MUX2X1 U10085 ( .B(n11810), .A(n11811), .S(n12602), .Y(n11809) );
  MUX2X1 U10086 ( .B(n11813), .A(n11814), .S(n12573), .Y(n11812) );
  MUX2X1 U10087 ( .B(n11816), .A(n11817), .S(n12602), .Y(n11815) );
  MUX2X1 U10088 ( .B(n11819), .A(n11820), .S(n12602), .Y(n11818) );
  MUX2X1 U10089 ( .B(n11822), .A(n11823), .S(n12602), .Y(n11821) );
  MUX2X1 U10090 ( .B(n11825), .A(n11826), .S(n12602), .Y(n11824) );
  MUX2X1 U10091 ( .B(n11828), .A(n11829), .S(n12573), .Y(n11827) );
  MUX2X1 U10092 ( .B(n11831), .A(n11832), .S(n12602), .Y(n11830) );
  MUX2X1 U10093 ( .B(n11834), .A(n11835), .S(n12602), .Y(n11833) );
  MUX2X1 U10094 ( .B(n11837), .A(n11838), .S(n12602), .Y(n11836) );
  MUX2X1 U10095 ( .B(n11840), .A(n11841), .S(n12602), .Y(n11839) );
  MUX2X1 U10096 ( .B(n11843), .A(n11844), .S(n12573), .Y(n11842) );
  MUX2X1 U10097 ( .B(n11846), .A(n11847), .S(n12603), .Y(n11845) );
  MUX2X1 U10098 ( .B(n11849), .A(n11850), .S(n12603), .Y(n11848) );
  MUX2X1 U10099 ( .B(n11852), .A(n11853), .S(n12603), .Y(n11851) );
  MUX2X1 U10100 ( .B(n11855), .A(n11856), .S(n12603), .Y(n11854) );
  MUX2X1 U10101 ( .B(n11858), .A(n11859), .S(n12573), .Y(n11857) );
  MUX2X1 U10102 ( .B(n11861), .A(n11862), .S(n12562), .Y(n11860) );
  MUX2X1 U10103 ( .B(n11864), .A(n11865), .S(n12603), .Y(n11863) );
  MUX2X1 U10104 ( .B(n11867), .A(n11868), .S(n12603), .Y(n11866) );
  MUX2X1 U10105 ( .B(n11870), .A(n11871), .S(n12603), .Y(n11869) );
  MUX2X1 U10106 ( .B(n11873), .A(n11874), .S(n12603), .Y(n11872) );
  MUX2X1 U10107 ( .B(n11876), .A(n11877), .S(n12573), .Y(n11875) );
  MUX2X1 U10108 ( .B(n11879), .A(n11880), .S(n12603), .Y(n11878) );
  MUX2X1 U10109 ( .B(n11882), .A(n11883), .S(n12603), .Y(n11881) );
  MUX2X1 U10110 ( .B(n11885), .A(n11886), .S(n12603), .Y(n11884) );
  MUX2X1 U10111 ( .B(n11888), .A(n11889), .S(n12603), .Y(n11887) );
  MUX2X1 U10112 ( .B(n11891), .A(n11892), .S(n12573), .Y(n11890) );
  MUX2X1 U10113 ( .B(n11894), .A(n11895), .S(n12604), .Y(n11893) );
  MUX2X1 U10114 ( .B(n11897), .A(n11898), .S(n12604), .Y(n11896) );
  MUX2X1 U10115 ( .B(n11900), .A(n11901), .S(n12604), .Y(n11899) );
  MUX2X1 U10116 ( .B(n11903), .A(n11904), .S(n12604), .Y(n11902) );
  MUX2X1 U10117 ( .B(n11906), .A(n11907), .S(n12573), .Y(n11905) );
  MUX2X1 U10118 ( .B(n11909), .A(n11910), .S(n12604), .Y(n11908) );
  MUX2X1 U10119 ( .B(n11912), .A(n11913), .S(n12604), .Y(n11911) );
  MUX2X1 U10120 ( .B(n11915), .A(n11916), .S(n12604), .Y(n11914) );
  MUX2X1 U10121 ( .B(n11918), .A(n11919), .S(n12604), .Y(n11917) );
  MUX2X1 U10122 ( .B(n11921), .A(n11922), .S(n12573), .Y(n11920) );
  MUX2X1 U10123 ( .B(n11924), .A(n11925), .S(n12563), .Y(n11923) );
  MUX2X1 U10124 ( .B(n11927), .A(n11928), .S(n12604), .Y(n11926) );
  MUX2X1 U10125 ( .B(n11930), .A(n11931), .S(n12604), .Y(n11929) );
  MUX2X1 U10126 ( .B(n11933), .A(n11934), .S(n12604), .Y(n11932) );
  MUX2X1 U10127 ( .B(n11936), .A(n11937), .S(n12604), .Y(n11935) );
  MUX2X1 U10128 ( .B(n11939), .A(n11940), .S(n12573), .Y(n11938) );
  MUX2X1 U10129 ( .B(n11942), .A(n11943), .S(n12605), .Y(n11941) );
  MUX2X1 U10130 ( .B(n11945), .A(n11946), .S(n12605), .Y(n11944) );
  MUX2X1 U10131 ( .B(n11948), .A(n11949), .S(n12605), .Y(n11947) );
  MUX2X1 U10132 ( .B(n11951), .A(n11952), .S(n12605), .Y(n11950) );
  MUX2X1 U10133 ( .B(n11954), .A(n11955), .S(n12573), .Y(n11953) );
  MUX2X1 U10134 ( .B(n11957), .A(n11958), .S(n12605), .Y(n11956) );
  MUX2X1 U10135 ( .B(n11960), .A(n11961), .S(n12605), .Y(n11959) );
  MUX2X1 U10136 ( .B(n11963), .A(n11964), .S(n12605), .Y(n11962) );
  MUX2X1 U10137 ( .B(n11966), .A(n11967), .S(n12605), .Y(n11965) );
  MUX2X1 U10138 ( .B(n11969), .A(n11970), .S(n12573), .Y(n11968) );
  MUX2X1 U10139 ( .B(n11972), .A(n11973), .S(n12605), .Y(n11971) );
  MUX2X1 U10140 ( .B(n11975), .A(n11976), .S(n12605), .Y(n11974) );
  MUX2X1 U10141 ( .B(n11978), .A(n11979), .S(n12605), .Y(n11977) );
  MUX2X1 U10142 ( .B(n11981), .A(n11982), .S(n12605), .Y(n11980) );
  MUX2X1 U10143 ( .B(n11984), .A(n11985), .S(n12573), .Y(n11983) );
  MUX2X1 U10144 ( .B(n11987), .A(n11988), .S(n12562), .Y(n11986) );
  MUX2X1 U10145 ( .B(n11990), .A(n11991), .S(n12606), .Y(n11989) );
  MUX2X1 U10146 ( .B(n11993), .A(n11994), .S(n12606), .Y(n11992) );
  MUX2X1 U10147 ( .B(n11996), .A(n11997), .S(n12606), .Y(n11995) );
  MUX2X1 U10148 ( .B(n11999), .A(n12000), .S(n12606), .Y(n11998) );
  MUX2X1 U10149 ( .B(n12002), .A(n12003), .S(n12571), .Y(n12001) );
  MUX2X1 U10150 ( .B(n12005), .A(n12006), .S(n12606), .Y(n12004) );
  MUX2X1 U10151 ( .B(n12008), .A(n12009), .S(n12606), .Y(n12007) );
  MUX2X1 U10152 ( .B(n12011), .A(n12012), .S(n12606), .Y(n12010) );
  MUX2X1 U10153 ( .B(n12014), .A(n12015), .S(n12606), .Y(n12013) );
  MUX2X1 U10154 ( .B(n12017), .A(n12018), .S(n12571), .Y(n12016) );
  MUX2X1 U10155 ( .B(n12020), .A(n12021), .S(n12606), .Y(n12019) );
  MUX2X1 U10156 ( .B(n12023), .A(n12024), .S(n12606), .Y(n12022) );
  MUX2X1 U10157 ( .B(n12026), .A(n12027), .S(n12606), .Y(n12025) );
  MUX2X1 U10158 ( .B(n12029), .A(n12030), .S(n12606), .Y(n12028) );
  MUX2X1 U10159 ( .B(n12032), .A(n12033), .S(n12571), .Y(n12031) );
  MUX2X1 U10160 ( .B(n12035), .A(n12036), .S(n12607), .Y(n12034) );
  MUX2X1 U10161 ( .B(n12038), .A(n12039), .S(n12607), .Y(n12037) );
  MUX2X1 U10162 ( .B(n12041), .A(n12042), .S(n12607), .Y(n12040) );
  MUX2X1 U10163 ( .B(n12044), .A(n12045), .S(n12607), .Y(n12043) );
  MUX2X1 U10164 ( .B(n12047), .A(n12048), .S(n12571), .Y(n12046) );
  MUX2X1 U10165 ( .B(n12050), .A(n12051), .S(n12562), .Y(n12049) );
  MUX2X1 U10166 ( .B(n12052), .A(n12053), .S(mem_access_addr[7]), .Y(
        mem_read_data[13]) );
  MUX2X1 U10167 ( .B(n12055), .A(n12056), .S(n12607), .Y(n12054) );
  MUX2X1 U10168 ( .B(n12058), .A(n12059), .S(n12607), .Y(n12057) );
  MUX2X1 U10169 ( .B(n12061), .A(n12062), .S(n12607), .Y(n12060) );
  MUX2X1 U10170 ( .B(n12064), .A(n12065), .S(n12607), .Y(n12063) );
  MUX2X1 U10171 ( .B(n12067), .A(n12068), .S(n12571), .Y(n12066) );
  MUX2X1 U10172 ( .B(n12070), .A(n12071), .S(n12607), .Y(n12069) );
  MUX2X1 U10173 ( .B(n12073), .A(n12074), .S(n12607), .Y(n12072) );
  MUX2X1 U10174 ( .B(n12076), .A(n12077), .S(n12607), .Y(n12075) );
  MUX2X1 U10175 ( .B(n12079), .A(n12080), .S(n12607), .Y(n12078) );
  MUX2X1 U10176 ( .B(n12082), .A(n12083), .S(n12571), .Y(n12081) );
  MUX2X1 U10177 ( .B(n12085), .A(n12086), .S(n12608), .Y(n12084) );
  MUX2X1 U10178 ( .B(n12088), .A(n12089), .S(n12608), .Y(n12087) );
  MUX2X1 U10179 ( .B(n12091), .A(n12092), .S(n12608), .Y(n12090) );
  MUX2X1 U10180 ( .B(n12094), .A(n12095), .S(n12608), .Y(n12093) );
  MUX2X1 U10181 ( .B(n12097), .A(n12098), .S(n12571), .Y(n12096) );
  MUX2X1 U10182 ( .B(n12100), .A(n12101), .S(n12608), .Y(n12099) );
  MUX2X1 U10183 ( .B(n12103), .A(n12104), .S(n12608), .Y(n12102) );
  MUX2X1 U10184 ( .B(n12106), .A(n12107), .S(n12608), .Y(n12105) );
  MUX2X1 U10185 ( .B(n12109), .A(n12110), .S(n12608), .Y(n12108) );
  MUX2X1 U10186 ( .B(n12112), .A(n12113), .S(n12571), .Y(n12111) );
  MUX2X1 U10187 ( .B(n12115), .A(n12116), .S(n12562), .Y(n12114) );
  MUX2X1 U10188 ( .B(n12118), .A(n12119), .S(n12608), .Y(n12117) );
  MUX2X1 U10189 ( .B(n12121), .A(n12122), .S(n12608), .Y(n12120) );
  MUX2X1 U10190 ( .B(n12124), .A(n12125), .S(n12608), .Y(n12123) );
  MUX2X1 U10191 ( .B(n12127), .A(n12128), .S(n12608), .Y(n12126) );
  MUX2X1 U10192 ( .B(n12130), .A(n12131), .S(n12571), .Y(n12129) );
  MUX2X1 U10193 ( .B(n12133), .A(n12134), .S(n12609), .Y(n12132) );
  MUX2X1 U10194 ( .B(n12136), .A(n12137), .S(n12609), .Y(n12135) );
  MUX2X1 U10195 ( .B(n12139), .A(n12140), .S(n12609), .Y(n12138) );
  MUX2X1 U10196 ( .B(n12142), .A(n12143), .S(n12609), .Y(n12141) );
  MUX2X1 U10197 ( .B(n12145), .A(n12146), .S(n12571), .Y(n12144) );
  MUX2X1 U10198 ( .B(n12148), .A(n12149), .S(n12609), .Y(n12147) );
  MUX2X1 U10199 ( .B(n12151), .A(n12152), .S(n12609), .Y(n12150) );
  MUX2X1 U10200 ( .B(n12154), .A(n12155), .S(n12609), .Y(n12153) );
  MUX2X1 U10201 ( .B(n12157), .A(n12158), .S(n12609), .Y(n12156) );
  MUX2X1 U10202 ( .B(n12160), .A(n12161), .S(n12571), .Y(n12159) );
  MUX2X1 U10203 ( .B(n12163), .A(n12164), .S(n12609), .Y(n12162) );
  MUX2X1 U10204 ( .B(n12166), .A(n12167), .S(n12609), .Y(n12165) );
  MUX2X1 U10205 ( .B(n12169), .A(n12170), .S(n12609), .Y(n12168) );
  MUX2X1 U10206 ( .B(n12172), .A(n12173), .S(n12609), .Y(n12171) );
  MUX2X1 U10207 ( .B(n12175), .A(n12176), .S(n12571), .Y(n12174) );
  MUX2X1 U10208 ( .B(n12178), .A(n12179), .S(n12563), .Y(n12177) );
  MUX2X1 U10209 ( .B(n12181), .A(n12182), .S(n12610), .Y(n12180) );
  MUX2X1 U10210 ( .B(n12184), .A(n12185), .S(n12610), .Y(n12183) );
  MUX2X1 U10211 ( .B(n12187), .A(n12188), .S(n12610), .Y(n12186) );
  MUX2X1 U10212 ( .B(n12190), .A(n12191), .S(n12610), .Y(n12189) );
  MUX2X1 U10213 ( .B(n12193), .A(n12194), .S(n12572), .Y(n12192) );
  MUX2X1 U10214 ( .B(n12196), .A(n12197), .S(n12610), .Y(n12195) );
  MUX2X1 U10215 ( .B(n12199), .A(n12200), .S(n12610), .Y(n12198) );
  MUX2X1 U10216 ( .B(n12202), .A(n12203), .S(n12610), .Y(n12201) );
  MUX2X1 U10217 ( .B(n12205), .A(n12206), .S(n12610), .Y(n12204) );
  MUX2X1 U10218 ( .B(n12208), .A(n12209), .S(n12572), .Y(n12207) );
  MUX2X1 U10219 ( .B(n12211), .A(n12212), .S(n12610), .Y(n12210) );
  MUX2X1 U10220 ( .B(n12214), .A(n12215), .S(n12610), .Y(n12213) );
  MUX2X1 U10221 ( .B(n12217), .A(n12218), .S(n12610), .Y(n12216) );
  MUX2X1 U10222 ( .B(n12220), .A(n12221), .S(n12610), .Y(n12219) );
  MUX2X1 U10223 ( .B(n12223), .A(n12224), .S(n12572), .Y(n12222) );
  MUX2X1 U10224 ( .B(n12226), .A(n12227), .S(n12611), .Y(n12225) );
  MUX2X1 U10225 ( .B(n12229), .A(n12230), .S(n12611), .Y(n12228) );
  MUX2X1 U10226 ( .B(n12232), .A(n12233), .S(n12611), .Y(n12231) );
  MUX2X1 U10227 ( .B(n12235), .A(n12236), .S(n12611), .Y(n12234) );
  MUX2X1 U10228 ( .B(n12238), .A(n12239), .S(n12572), .Y(n12237) );
  MUX2X1 U10229 ( .B(n12241), .A(n12242), .S(n12562), .Y(n12240) );
  MUX2X1 U10230 ( .B(n12244), .A(n12245), .S(n12611), .Y(n12243) );
  MUX2X1 U10231 ( .B(n12247), .A(n12248), .S(n12611), .Y(n12246) );
  MUX2X1 U10232 ( .B(n12250), .A(n12251), .S(n12611), .Y(n12249) );
  MUX2X1 U10233 ( .B(n12253), .A(n12254), .S(n12611), .Y(n12252) );
  MUX2X1 U10234 ( .B(n12256), .A(n12257), .S(n12572), .Y(n12255) );
  MUX2X1 U10235 ( .B(n12259), .A(n12260), .S(n12611), .Y(n12258) );
  MUX2X1 U10236 ( .B(n12262), .A(n12263), .S(n12611), .Y(n12261) );
  MUX2X1 U10237 ( .B(n12265), .A(n12266), .S(n12611), .Y(n12264) );
  MUX2X1 U10238 ( .B(n12268), .A(n12269), .S(n12611), .Y(n12267) );
  MUX2X1 U10239 ( .B(n12271), .A(n12272), .S(n12572), .Y(n12270) );
  MUX2X1 U10240 ( .B(n12274), .A(n12275), .S(n12612), .Y(n12273) );
  MUX2X1 U10241 ( .B(n12277), .A(n12278), .S(n12612), .Y(n12276) );
  MUX2X1 U10242 ( .B(n12280), .A(n12281), .S(n12612), .Y(n12279) );
  MUX2X1 U10243 ( .B(n12283), .A(n12284), .S(n12612), .Y(n12282) );
  MUX2X1 U10244 ( .B(n12286), .A(n12287), .S(n12572), .Y(n12285) );
  MUX2X1 U10245 ( .B(n12289), .A(n12290), .S(n12612), .Y(n12288) );
  MUX2X1 U10246 ( .B(n12292), .A(n12293), .S(n12612), .Y(n12291) );
  MUX2X1 U10247 ( .B(n12295), .A(n12296), .S(n12612), .Y(n12294) );
  MUX2X1 U10248 ( .B(n12298), .A(n12299), .S(n12612), .Y(n12297) );
  MUX2X1 U10249 ( .B(n12301), .A(n12302), .S(n12572), .Y(n12300) );
  MUX2X1 U10250 ( .B(n12304), .A(n12305), .S(n12562), .Y(n12303) );
  MUX2X1 U10251 ( .B(n12306), .A(n12307), .S(mem_access_addr[7]), .Y(
        mem_read_data[14]) );
  MUX2X1 U10252 ( .B(n12309), .A(n12310), .S(n12612), .Y(n12308) );
  MUX2X1 U10253 ( .B(n12312), .A(n12313), .S(n12612), .Y(n12311) );
  MUX2X1 U10254 ( .B(n12315), .A(n12316), .S(n12612), .Y(n12314) );
  MUX2X1 U10255 ( .B(n12318), .A(n12319), .S(n12612), .Y(n12317) );
  MUX2X1 U10256 ( .B(n12321), .A(n12322), .S(n12572), .Y(n12320) );
  MUX2X1 U10257 ( .B(n12324), .A(n12325), .S(n12613), .Y(n12323) );
  MUX2X1 U10258 ( .B(n12327), .A(n12328), .S(n12613), .Y(n12326) );
  MUX2X1 U10259 ( .B(n12330), .A(n12331), .S(n12613), .Y(n12329) );
  MUX2X1 U10260 ( .B(n12333), .A(n12334), .S(n12613), .Y(n12332) );
  MUX2X1 U10261 ( .B(n12336), .A(n12337), .S(n12572), .Y(n12335) );
  MUX2X1 U10262 ( .B(n12339), .A(n12340), .S(n12613), .Y(n12338) );
  MUX2X1 U10263 ( .B(n12342), .A(n12343), .S(n12613), .Y(n12341) );
  MUX2X1 U10264 ( .B(n12345), .A(n12346), .S(n12613), .Y(n12344) );
  MUX2X1 U10265 ( .B(n12348), .A(n12349), .S(n12613), .Y(n12347) );
  MUX2X1 U10266 ( .B(n12351), .A(n12352), .S(n12572), .Y(n12350) );
  MUX2X1 U10267 ( .B(n12354), .A(n12355), .S(n12613), .Y(n12353) );
  MUX2X1 U10268 ( .B(n12357), .A(n12358), .S(n12613), .Y(n12356) );
  MUX2X1 U10269 ( .B(n12360), .A(n12361), .S(n12613), .Y(n12359) );
  MUX2X1 U10270 ( .B(n12363), .A(n12364), .S(n12613), .Y(n12362) );
  MUX2X1 U10271 ( .B(n12366), .A(n12367), .S(n12572), .Y(n12365) );
  MUX2X1 U10272 ( .B(n12369), .A(n12370), .S(n12562), .Y(n12368) );
  MUX2X1 U10273 ( .B(n12372), .A(n12373), .S(n12614), .Y(n12371) );
  MUX2X1 U10274 ( .B(n12375), .A(n12376), .S(n12614), .Y(n12374) );
  MUX2X1 U10275 ( .B(n12378), .A(n12379), .S(n12614), .Y(n12377) );
  MUX2X1 U10276 ( .B(n12381), .A(n12382), .S(n12614), .Y(n12380) );
  MUX2X1 U10277 ( .B(n12384), .A(n12385), .S(n12573), .Y(n12383) );
  MUX2X1 U10278 ( .B(n12387), .A(n12388), .S(n12614), .Y(n12386) );
  MUX2X1 U10279 ( .B(n12390), .A(n12391), .S(n12614), .Y(n12389) );
  MUX2X1 U10280 ( .B(n12393), .A(n12394), .S(n12614), .Y(n12392) );
  MUX2X1 U10281 ( .B(n12396), .A(n12397), .S(n12614), .Y(n12395) );
  MUX2X1 U10282 ( .B(n12399), .A(n12400), .S(n12573), .Y(n12398) );
  MUX2X1 U10283 ( .B(n12402), .A(n12403), .S(n12614), .Y(n12401) );
  MUX2X1 U10284 ( .B(n12405), .A(n12406), .S(n12614), .Y(n12404) );
  MUX2X1 U10285 ( .B(n12408), .A(n12409), .S(n12614), .Y(n12407) );
  MUX2X1 U10286 ( .B(n12411), .A(n12412), .S(n12614), .Y(n12410) );
  MUX2X1 U10287 ( .B(n12414), .A(n12415), .S(n12573), .Y(n12413) );
  MUX2X1 U10288 ( .B(n12417), .A(n12418), .S(n12615), .Y(n12416) );
  MUX2X1 U10289 ( .B(n12420), .A(n12421), .S(n12615), .Y(n12419) );
  MUX2X1 U10290 ( .B(n12423), .A(n12424), .S(n12615), .Y(n12422) );
  MUX2X1 U10291 ( .B(n12426), .A(n12427), .S(n12615), .Y(n12425) );
  MUX2X1 U10292 ( .B(n12429), .A(n12430), .S(n12573), .Y(n12428) );
  MUX2X1 U10293 ( .B(n12432), .A(n12433), .S(n12562), .Y(n12431) );
  MUX2X1 U10294 ( .B(n12435), .A(n12436), .S(n12615), .Y(n12434) );
  MUX2X1 U10295 ( .B(n12438), .A(n12439), .S(n12615), .Y(n12437) );
  MUX2X1 U10296 ( .B(n12441), .A(n12442), .S(n12615), .Y(n12440) );
  MUX2X1 U10297 ( .B(n12444), .A(n12445), .S(n12615), .Y(n12443) );
  MUX2X1 U10298 ( .B(n12447), .A(n12448), .S(n12573), .Y(n12446) );
  MUX2X1 U10299 ( .B(n12450), .A(n12451), .S(n12615), .Y(n12449) );
  MUX2X1 U10300 ( .B(n12453), .A(n12454), .S(n12615), .Y(n12452) );
  MUX2X1 U10301 ( .B(n12456), .A(n12457), .S(n12615), .Y(n12455) );
  MUX2X1 U10302 ( .B(n12459), .A(n12460), .S(n12615), .Y(n12458) );
  MUX2X1 U10303 ( .B(n12462), .A(n12463), .S(n12573), .Y(n12461) );
  MUX2X1 U10304 ( .B(n12465), .A(n12466), .S(n12616), .Y(n12464) );
  MUX2X1 U10305 ( .B(n12468), .A(n12469), .S(n12616), .Y(n12467) );
  MUX2X1 U10306 ( .B(n12471), .A(n12472), .S(n12616), .Y(n12470) );
  MUX2X1 U10307 ( .B(n12474), .A(n12475), .S(n12616), .Y(n12473) );
  MUX2X1 U10308 ( .B(n12477), .A(n12478), .S(n12573), .Y(n12476) );
  MUX2X1 U10309 ( .B(n12480), .A(n12481), .S(n12616), .Y(n12479) );
  MUX2X1 U10310 ( .B(n12483), .A(n12484), .S(n12616), .Y(n12482) );
  MUX2X1 U10311 ( .B(n12486), .A(n12487), .S(n12616), .Y(n12485) );
  MUX2X1 U10312 ( .B(n12489), .A(n12490), .S(n12616), .Y(n12488) );
  MUX2X1 U10313 ( .B(n12492), .A(n12493), .S(n12573), .Y(n12491) );
  MUX2X1 U10314 ( .B(n12495), .A(n12496), .S(n12562), .Y(n12494) );
  MUX2X1 U10315 ( .B(n12498), .A(n12499), .S(n12616), .Y(n12497) );
  MUX2X1 U10316 ( .B(n12501), .A(n12502), .S(n12616), .Y(n12500) );
  MUX2X1 U10317 ( .B(n12504), .A(n12505), .S(n12616), .Y(n12503) );
  MUX2X1 U10318 ( .B(n12507), .A(n12508), .S(n12616), .Y(n12506) );
  MUX2X1 U10319 ( .B(n12510), .A(n12511), .S(n12573), .Y(n12509) );
  MUX2X1 U10320 ( .B(n12513), .A(n12514), .S(n12617), .Y(n12512) );
  MUX2X1 U10321 ( .B(n12516), .A(n12517), .S(n12617), .Y(n12515) );
  MUX2X1 U10322 ( .B(n12519), .A(n12520), .S(n12617), .Y(n12518) );
  MUX2X1 U10323 ( .B(n12522), .A(n12523), .S(n12617), .Y(n12521) );
  MUX2X1 U10324 ( .B(n12525), .A(n12526), .S(n12573), .Y(n12524) );
  MUX2X1 U10325 ( .B(n12528), .A(n12529), .S(n12617), .Y(n12527) );
  MUX2X1 U10326 ( .B(n12531), .A(n12532), .S(n12617), .Y(n12530) );
  MUX2X1 U10327 ( .B(n12534), .A(n12535), .S(n12617), .Y(n12533) );
  MUX2X1 U10328 ( .B(n12537), .A(n12538), .S(n12617), .Y(n12536) );
  MUX2X1 U10329 ( .B(n12540), .A(n12541), .S(n12573), .Y(n12539) );
  MUX2X1 U10330 ( .B(n12543), .A(n12544), .S(n12617), .Y(n12542) );
  MUX2X1 U10331 ( .B(n12546), .A(n12547), .S(n12617), .Y(n12545) );
  MUX2X1 U10332 ( .B(n12549), .A(n12550), .S(n12617), .Y(n12548) );
  MUX2X1 U10333 ( .B(n12552), .A(n12553), .S(n12617), .Y(n12551) );
  MUX2X1 U10334 ( .B(n12555), .A(n12556), .S(n12573), .Y(n12554) );
  MUX2X1 U10335 ( .B(n12558), .A(n12559), .S(n12563), .Y(n12557) );
  MUX2X1 U10336 ( .B(n12560), .A(n12561), .S(mem_access_addr[7]), .Y(
        mem_read_data[15]) );
  MUX2X1 U10337 ( .B(ram[4064]), .A(ram[4080]), .S(n12639), .Y(n3865) );
  MUX2X1 U10338 ( .B(ram[4032]), .A(ram[4048]), .S(n12639), .Y(n3848) );
  MUX2X1 U10339 ( .B(ram[4000]), .A(ram[4016]), .S(n12639), .Y(n3917) );
  MUX2X1 U10340 ( .B(ram[3968]), .A(ram[3984]), .S(n12639), .Y(n3900) );
  MUX2X1 U10341 ( .B(n3883), .A(n3831), .S(n12589), .Y(n4070) );
  MUX2X1 U10342 ( .B(ram[3936]), .A(ram[3952]), .S(n12639), .Y(n3968) );
  MUX2X1 U10343 ( .B(ram[3904]), .A(ram[3920]), .S(n12639), .Y(n3951) );
  MUX2X1 U10344 ( .B(ram[3872]), .A(ram[3888]), .S(n12639), .Y(n4019) );
  MUX2X1 U10345 ( .B(ram[3840]), .A(ram[3856]), .S(n12639), .Y(n4002) );
  MUX2X1 U10346 ( .B(n3985), .A(n3934), .S(mem_access_addr[2]), .Y(n4053) );
  MUX2X1 U10347 ( .B(ram[3808]), .A(ram[3824]), .S(n12640), .Y(n4121) );
  MUX2X1 U10348 ( .B(ram[3776]), .A(ram[3792]), .S(n12640), .Y(n4104) );
  MUX2X1 U10349 ( .B(ram[3744]), .A(ram[3760]), .S(n12640), .Y(n4175) );
  MUX2X1 U10350 ( .B(ram[3712]), .A(ram[3728]), .S(n12640), .Y(n4156) );
  MUX2X1 U10351 ( .B(n4138), .A(n4087), .S(n12586), .Y(n4333) );
  MUX2X1 U10352 ( .B(ram[3680]), .A(ram[3696]), .S(n12640), .Y(n4229) );
  MUX2X1 U10353 ( .B(ram[3648]), .A(ram[3664]), .S(n12640), .Y(n4211) );
  MUX2X1 U10354 ( .B(ram[3616]), .A(ram[3632]), .S(n12640), .Y(n4281) );
  MUX2X1 U10355 ( .B(ram[3584]), .A(ram[3600]), .S(n12640), .Y(n4264) );
  MUX2X1 U10356 ( .B(n4247), .A(n4193), .S(n12579), .Y(n4316) );
  MUX2X1 U10357 ( .B(n4298), .A(n4036), .S(n12564), .Y(n8560) );
  MUX2X1 U10358 ( .B(ram[3552]), .A(ram[3568]), .S(n12640), .Y(n4385) );
  MUX2X1 U10359 ( .B(ram[3520]), .A(ram[3536]), .S(n12640), .Y(n4367) );
  MUX2X1 U10360 ( .B(ram[3488]), .A(ram[3504]), .S(n12640), .Y(n8533) );
  MUX2X1 U10361 ( .B(ram[3456]), .A(ram[3472]), .S(n12640), .Y(n4419) );
  MUX2X1 U10362 ( .B(n4402), .A(n4350), .S(mem_access_addr[2]), .Y(n8542) );
  MUX2X1 U10363 ( .B(ram[3424]), .A(ram[3440]), .S(n12641), .Y(n8536) );
  MUX2X1 U10364 ( .B(ram[3392]), .A(ram[3408]), .S(n12641), .Y(n8535) );
  MUX2X1 U10365 ( .B(ram[3360]), .A(ram[3376]), .S(n12641), .Y(n8539) );
  MUX2X1 U10366 ( .B(ram[3328]), .A(ram[3344]), .S(n12641), .Y(n8538) );
  MUX2X1 U10367 ( .B(n8537), .A(n8534), .S(mem_access_addr[2]), .Y(n8541) );
  MUX2X1 U10368 ( .B(ram[3296]), .A(ram[3312]), .S(n12641), .Y(n8545) );
  MUX2X1 U10369 ( .B(ram[3264]), .A(ram[3280]), .S(n12641), .Y(n8544) );
  MUX2X1 U10370 ( .B(ram[3232]), .A(ram[3248]), .S(n12641), .Y(n8548) );
  MUX2X1 U10371 ( .B(ram[3200]), .A(ram[3216]), .S(n12641), .Y(n8547) );
  MUX2X1 U10372 ( .B(n8546), .A(n8543), .S(n12587), .Y(n8557) );
  MUX2X1 U10373 ( .B(ram[3168]), .A(ram[3184]), .S(n12641), .Y(n8551) );
  MUX2X1 U10374 ( .B(ram[3136]), .A(ram[3152]), .S(n12641), .Y(n8550) );
  MUX2X1 U10375 ( .B(ram[3104]), .A(ram[3120]), .S(n12641), .Y(n8554) );
  MUX2X1 U10376 ( .B(ram[3072]), .A(ram[3088]), .S(n12641), .Y(n8553) );
  MUX2X1 U10377 ( .B(n8552), .A(n8549), .S(mem_access_addr[2]), .Y(n8556) );
  MUX2X1 U10378 ( .B(n8555), .A(n8540), .S(n12564), .Y(n8559) );
  MUX2X1 U10379 ( .B(ram[3040]), .A(ram[3056]), .S(n12642), .Y(n8563) );
  MUX2X1 U10380 ( .B(ram[3008]), .A(ram[3024]), .S(n12642), .Y(n8562) );
  MUX2X1 U10381 ( .B(ram[2976]), .A(ram[2992]), .S(n12642), .Y(n8566) );
  MUX2X1 U10382 ( .B(ram[2944]), .A(ram[2960]), .S(n12642), .Y(n8565) );
  MUX2X1 U10383 ( .B(n8564), .A(n8561), .S(n12579), .Y(n8575) );
  MUX2X1 U10384 ( .B(ram[2912]), .A(ram[2928]), .S(n12642), .Y(n8569) );
  MUX2X1 U10385 ( .B(ram[2880]), .A(ram[2896]), .S(n12642), .Y(n8568) );
  MUX2X1 U10386 ( .B(ram[2848]), .A(ram[2864]), .S(n12642), .Y(n8572) );
  MUX2X1 U10387 ( .B(ram[2816]), .A(ram[2832]), .S(n12642), .Y(n8571) );
  MUX2X1 U10388 ( .B(n8570), .A(n8567), .S(n12585), .Y(n8574) );
  MUX2X1 U10389 ( .B(ram[2784]), .A(ram[2800]), .S(n12642), .Y(n8578) );
  MUX2X1 U10390 ( .B(ram[2752]), .A(ram[2768]), .S(n12642), .Y(n8577) );
  MUX2X1 U10391 ( .B(ram[2720]), .A(ram[2736]), .S(n12642), .Y(n8581) );
  MUX2X1 U10392 ( .B(ram[2688]), .A(ram[2704]), .S(n12642), .Y(n8580) );
  MUX2X1 U10393 ( .B(n8579), .A(n8576), .S(n12578), .Y(n8590) );
  MUX2X1 U10394 ( .B(ram[2656]), .A(ram[2672]), .S(n12643), .Y(n8584) );
  MUX2X1 U10395 ( .B(ram[2624]), .A(ram[2640]), .S(n12643), .Y(n8583) );
  MUX2X1 U10396 ( .B(ram[2592]), .A(ram[2608]), .S(n12643), .Y(n8587) );
  MUX2X1 U10397 ( .B(ram[2560]), .A(ram[2576]), .S(n12643), .Y(n8586) );
  MUX2X1 U10398 ( .B(n8585), .A(n8582), .S(n12582), .Y(n8589) );
  MUX2X1 U10399 ( .B(n8588), .A(n8573), .S(n12564), .Y(n8623) );
  MUX2X1 U10400 ( .B(ram[2528]), .A(ram[2544]), .S(n12643), .Y(n8593) );
  MUX2X1 U10401 ( .B(ram[2496]), .A(ram[2512]), .S(n12643), .Y(n8592) );
  MUX2X1 U10402 ( .B(ram[2464]), .A(ram[2480]), .S(n12643), .Y(n8596) );
  MUX2X1 U10403 ( .B(ram[2432]), .A(ram[2448]), .S(n12643), .Y(n8595) );
  MUX2X1 U10404 ( .B(n8594), .A(n8591), .S(n12583), .Y(n8605) );
  MUX2X1 U10405 ( .B(ram[2400]), .A(ram[2416]), .S(n12643), .Y(n8599) );
  MUX2X1 U10406 ( .B(ram[2368]), .A(ram[2384]), .S(n12643), .Y(n8598) );
  MUX2X1 U10407 ( .B(ram[2336]), .A(ram[2352]), .S(n12643), .Y(n8602) );
  MUX2X1 U10408 ( .B(ram[2304]), .A(ram[2320]), .S(n12643), .Y(n8601) );
  MUX2X1 U10409 ( .B(n8600), .A(n8597), .S(n12579), .Y(n8604) );
  MUX2X1 U10410 ( .B(ram[2272]), .A(ram[2288]), .S(n12644), .Y(n8608) );
  MUX2X1 U10411 ( .B(ram[2240]), .A(ram[2256]), .S(n12644), .Y(n8607) );
  MUX2X1 U10412 ( .B(ram[2208]), .A(ram[2224]), .S(n12644), .Y(n8611) );
  MUX2X1 U10413 ( .B(ram[2176]), .A(ram[2192]), .S(n12644), .Y(n8610) );
  MUX2X1 U10414 ( .B(n8609), .A(n8606), .S(n12580), .Y(n8620) );
  MUX2X1 U10415 ( .B(ram[2144]), .A(ram[2160]), .S(n12644), .Y(n8614) );
  MUX2X1 U10416 ( .B(ram[2112]), .A(ram[2128]), .S(n12644), .Y(n8613) );
  MUX2X1 U10417 ( .B(ram[2080]), .A(ram[2096]), .S(n12644), .Y(n8617) );
  MUX2X1 U10418 ( .B(ram[2048]), .A(ram[2064]), .S(n12644), .Y(n8616) );
  MUX2X1 U10419 ( .B(n8615), .A(n8612), .S(n12575), .Y(n8619) );
  MUX2X1 U10420 ( .B(n8618), .A(n8603), .S(n12564), .Y(n8622) );
  MUX2X1 U10421 ( .B(n8621), .A(n8558), .S(mem_access_addr[6]), .Y(n8751) );
  MUX2X1 U10422 ( .B(ram[2016]), .A(ram[2032]), .S(n12644), .Y(n8626) );
  MUX2X1 U10423 ( .B(ram[1984]), .A(ram[2000]), .S(n12644), .Y(n8625) );
  MUX2X1 U10424 ( .B(ram[1952]), .A(ram[1968]), .S(n12644), .Y(n8629) );
  MUX2X1 U10425 ( .B(ram[1920]), .A(ram[1936]), .S(n12644), .Y(n8628) );
  MUX2X1 U10426 ( .B(n8627), .A(n8624), .S(n12577), .Y(n8638) );
  MUX2X1 U10427 ( .B(ram[1888]), .A(ram[1904]), .S(n12645), .Y(n8632) );
  MUX2X1 U10428 ( .B(ram[1856]), .A(ram[1872]), .S(n12645), .Y(n8631) );
  MUX2X1 U10429 ( .B(ram[1824]), .A(ram[1840]), .S(n12645), .Y(n8635) );
  MUX2X1 U10430 ( .B(ram[1792]), .A(ram[1808]), .S(n12645), .Y(n8634) );
  MUX2X1 U10431 ( .B(n8633), .A(n8630), .S(n12578), .Y(n8637) );
  MUX2X1 U10432 ( .B(ram[1760]), .A(ram[1776]), .S(n12645), .Y(n8641) );
  MUX2X1 U10433 ( .B(ram[1728]), .A(ram[1744]), .S(n12645), .Y(n8640) );
  MUX2X1 U10434 ( .B(ram[1696]), .A(ram[1712]), .S(n12645), .Y(n8644) );
  MUX2X1 U10435 ( .B(ram[1664]), .A(ram[1680]), .S(n12645), .Y(n8643) );
  MUX2X1 U10436 ( .B(n8642), .A(n8639), .S(n12586), .Y(n8653) );
  MUX2X1 U10437 ( .B(ram[1632]), .A(ram[1648]), .S(n12645), .Y(n8647) );
  MUX2X1 U10438 ( .B(ram[1600]), .A(ram[1616]), .S(n12645), .Y(n8646) );
  MUX2X1 U10439 ( .B(ram[1568]), .A(ram[1584]), .S(n12645), .Y(n8650) );
  MUX2X1 U10440 ( .B(ram[1536]), .A(ram[1552]), .S(n12645), .Y(n8649) );
  MUX2X1 U10441 ( .B(n8648), .A(n8645), .S(n12576), .Y(n8652) );
  MUX2X1 U10442 ( .B(n8651), .A(n8636), .S(n12564), .Y(n8686) );
  MUX2X1 U10443 ( .B(ram[1504]), .A(ram[1520]), .S(n12646), .Y(n8656) );
  MUX2X1 U10444 ( .B(ram[1472]), .A(ram[1488]), .S(n12646), .Y(n8655) );
  MUX2X1 U10445 ( .B(ram[1440]), .A(ram[1456]), .S(n12646), .Y(n8659) );
  MUX2X1 U10446 ( .B(ram[1408]), .A(ram[1424]), .S(n12646), .Y(n8658) );
  MUX2X1 U10447 ( .B(n8657), .A(n8654), .S(mem_access_addr[2]), .Y(n8668) );
  MUX2X1 U10448 ( .B(ram[1376]), .A(ram[1392]), .S(n12646), .Y(n8662) );
  MUX2X1 U10449 ( .B(ram[1344]), .A(ram[1360]), .S(n12646), .Y(n8661) );
  MUX2X1 U10450 ( .B(ram[1312]), .A(ram[1328]), .S(n12646), .Y(n8665) );
  MUX2X1 U10451 ( .B(ram[1280]), .A(ram[1296]), .S(n12646), .Y(n8664) );
  MUX2X1 U10452 ( .B(n8663), .A(n8660), .S(mem_access_addr[2]), .Y(n8667) );
  MUX2X1 U10453 ( .B(ram[1248]), .A(ram[1264]), .S(n12646), .Y(n8671) );
  MUX2X1 U10454 ( .B(ram[1216]), .A(ram[1232]), .S(n12646), .Y(n8670) );
  MUX2X1 U10455 ( .B(ram[1184]), .A(ram[1200]), .S(n12646), .Y(n8674) );
  MUX2X1 U10456 ( .B(ram[1152]), .A(ram[1168]), .S(n12646), .Y(n8673) );
  MUX2X1 U10457 ( .B(n8672), .A(n8669), .S(mem_access_addr[2]), .Y(n8683) );
  MUX2X1 U10458 ( .B(ram[1120]), .A(ram[1136]), .S(n12647), .Y(n8677) );
  MUX2X1 U10459 ( .B(ram[1088]), .A(ram[1104]), .S(n12647), .Y(n8676) );
  MUX2X1 U10460 ( .B(ram[1056]), .A(ram[1072]), .S(n12647), .Y(n8680) );
  MUX2X1 U10461 ( .B(ram[1024]), .A(ram[1040]), .S(n12647), .Y(n8679) );
  MUX2X1 U10462 ( .B(n8678), .A(n8675), .S(mem_access_addr[2]), .Y(n8682) );
  MUX2X1 U10463 ( .B(n8681), .A(n8666), .S(n12564), .Y(n8685) );
  MUX2X1 U10464 ( .B(ram[992]), .A(ram[1008]), .S(n12647), .Y(n8689) );
  MUX2X1 U10465 ( .B(ram[960]), .A(ram[976]), .S(n12647), .Y(n8688) );
  MUX2X1 U10466 ( .B(ram[928]), .A(ram[944]), .S(n12647), .Y(n8692) );
  MUX2X1 U10467 ( .B(ram[896]), .A(ram[912]), .S(n12647), .Y(n8691) );
  MUX2X1 U10468 ( .B(n8690), .A(n8687), .S(n12583), .Y(n8701) );
  MUX2X1 U10469 ( .B(ram[864]), .A(ram[880]), .S(n12647), .Y(n8695) );
  MUX2X1 U10470 ( .B(ram[832]), .A(ram[848]), .S(n12647), .Y(n8694) );
  MUX2X1 U10471 ( .B(ram[800]), .A(ram[816]), .S(n12647), .Y(n8698) );
  MUX2X1 U10472 ( .B(ram[768]), .A(ram[784]), .S(n12647), .Y(n8697) );
  MUX2X1 U10473 ( .B(n8696), .A(n8693), .S(mem_access_addr[2]), .Y(n8700) );
  MUX2X1 U10474 ( .B(ram[736]), .A(ram[752]), .S(n12669), .Y(n8704) );
  MUX2X1 U10475 ( .B(ram[704]), .A(ram[720]), .S(n12663), .Y(n8703) );
  MUX2X1 U10476 ( .B(ram[672]), .A(ram[688]), .S(n12625), .Y(n8707) );
  MUX2X1 U10477 ( .B(ram[640]), .A(ram[656]), .S(n12626), .Y(n8706) );
  MUX2X1 U10478 ( .B(n8705), .A(n8702), .S(n12589), .Y(n8716) );
  MUX2X1 U10479 ( .B(ram[608]), .A(ram[624]), .S(n12635), .Y(n8710) );
  MUX2X1 U10480 ( .B(ram[576]), .A(ram[592]), .S(n12645), .Y(n8709) );
  MUX2X1 U10481 ( .B(ram[544]), .A(ram[560]), .S(n12633), .Y(n8713) );
  MUX2X1 U10482 ( .B(ram[512]), .A(ram[528]), .S(n12671), .Y(n8712) );
  MUX2X1 U10483 ( .B(n8711), .A(n8708), .S(n12583), .Y(n8715) );
  MUX2X1 U10484 ( .B(n8714), .A(n8699), .S(n12564), .Y(n8749) );
  MUX2X1 U10485 ( .B(ram[480]), .A(ram[496]), .S(n12647), .Y(n8719) );
  MUX2X1 U10486 ( .B(ram[448]), .A(ram[464]), .S(n12682), .Y(n8718) );
  MUX2X1 U10487 ( .B(ram[416]), .A(ram[432]), .S(n12625), .Y(n8722) );
  MUX2X1 U10488 ( .B(ram[384]), .A(ram[400]), .S(n12650), .Y(n8721) );
  MUX2X1 U10489 ( .B(n8720), .A(n8717), .S(mem_access_addr[2]), .Y(n8731) );
  MUX2X1 U10490 ( .B(ram[352]), .A(ram[368]), .S(n12659), .Y(n8725) );
  MUX2X1 U10491 ( .B(ram[320]), .A(ram[336]), .S(n12639), .Y(n8724) );
  MUX2X1 U10492 ( .B(ram[288]), .A(ram[304]), .S(n12682), .Y(n8728) );
  MUX2X1 U10493 ( .B(ram[256]), .A(ram[272]), .S(n12628), .Y(n8727) );
  MUX2X1 U10494 ( .B(n8726), .A(n8723), .S(mem_access_addr[2]), .Y(n8730) );
  MUX2X1 U10495 ( .B(ram[224]), .A(ram[240]), .S(n12683), .Y(n8734) );
  MUX2X1 U10496 ( .B(ram[192]), .A(ram[208]), .S(n12675), .Y(n8733) );
  MUX2X1 U10497 ( .B(ram[160]), .A(ram[176]), .S(n12628), .Y(n8737) );
  MUX2X1 U10498 ( .B(ram[128]), .A(ram[144]), .S(n12647), .Y(n8736) );
  MUX2X1 U10499 ( .B(n8735), .A(n8732), .S(n12581), .Y(n8746) );
  MUX2X1 U10500 ( .B(ram[96]), .A(ram[112]), .S(n12656), .Y(n8740) );
  MUX2X1 U10501 ( .B(ram[64]), .A(ram[80]), .S(n12644), .Y(n8739) );
  MUX2X1 U10502 ( .B(ram[32]), .A(ram[48]), .S(n12641), .Y(n8743) );
  MUX2X1 U10503 ( .B(ram[0]), .A(ram[16]), .S(n12663), .Y(n8742) );
  MUX2X1 U10504 ( .B(n8741), .A(n8738), .S(mem_access_addr[2]), .Y(n8745) );
  MUX2X1 U10505 ( .B(n8744), .A(n8729), .S(n12564), .Y(n8748) );
  MUX2X1 U10506 ( .B(n8747), .A(n8684), .S(n1), .Y(n8750) );
  MUX2X1 U10507 ( .B(ram[4065]), .A(ram[4081]), .S(n12630), .Y(n8754) );
  MUX2X1 U10508 ( .B(ram[4033]), .A(ram[4049]), .S(n12642), .Y(n8753) );
  MUX2X1 U10509 ( .B(ram[4001]), .A(ram[4017]), .S(n12648), .Y(n8757) );
  MUX2X1 U10510 ( .B(ram[3969]), .A(ram[3985]), .S(n12650), .Y(n8756) );
  MUX2X1 U10511 ( .B(n8755), .A(n8752), .S(n12576), .Y(n8766) );
  MUX2X1 U10512 ( .B(ram[3937]), .A(ram[3953]), .S(n12626), .Y(n8760) );
  MUX2X1 U10513 ( .B(ram[3905]), .A(ram[3921]), .S(n12670), .Y(n8759) );
  MUX2X1 U10514 ( .B(ram[3873]), .A(ram[3889]), .S(n12666), .Y(n8763) );
  MUX2X1 U10515 ( .B(ram[3841]), .A(ram[3857]), .S(n12683), .Y(n8762) );
  MUX2X1 U10516 ( .B(n8761), .A(n8758), .S(n12585), .Y(n8765) );
  MUX2X1 U10517 ( .B(ram[3809]), .A(ram[3825]), .S(n12627), .Y(n8769) );
  MUX2X1 U10518 ( .B(ram[3777]), .A(ram[3793]), .S(n12647), .Y(n8768) );
  MUX2X1 U10519 ( .B(ram[3745]), .A(ram[3761]), .S(n12626), .Y(n8772) );
  MUX2X1 U10520 ( .B(ram[3713]), .A(ram[3729]), .S(n12639), .Y(n8771) );
  MUX2X1 U10521 ( .B(n8770), .A(n8767), .S(n12587), .Y(n8781) );
  MUX2X1 U10522 ( .B(ram[3681]), .A(ram[3697]), .S(n12660), .Y(n8775) );
  MUX2X1 U10523 ( .B(ram[3649]), .A(ram[3665]), .S(n12668), .Y(n8774) );
  MUX2X1 U10524 ( .B(ram[3617]), .A(ram[3633]), .S(n12680), .Y(n8778) );
  MUX2X1 U10525 ( .B(ram[3585]), .A(ram[3601]), .S(n12672), .Y(n8777) );
  MUX2X1 U10526 ( .B(n8776), .A(n8773), .S(n12583), .Y(n8780) );
  MUX2X1 U10527 ( .B(n8779), .A(n8764), .S(n12564), .Y(n8814) );
  MUX2X1 U10528 ( .B(ram[3553]), .A(ram[3569]), .S(n12675), .Y(n8784) );
  MUX2X1 U10529 ( .B(ram[3521]), .A(ram[3537]), .S(n12621), .Y(n8783) );
  MUX2X1 U10530 ( .B(ram[3489]), .A(ram[3505]), .S(n12680), .Y(n8787) );
  MUX2X1 U10531 ( .B(ram[3457]), .A(ram[3473]), .S(n12660), .Y(n8786) );
  MUX2X1 U10532 ( .B(n8785), .A(n8782), .S(n12584), .Y(n8796) );
  MUX2X1 U10533 ( .B(ram[3425]), .A(ram[3441]), .S(n12681), .Y(n8790) );
  MUX2X1 U10534 ( .B(ram[3393]), .A(ram[3409]), .S(n12670), .Y(n8789) );
  MUX2X1 U10535 ( .B(ram[3361]), .A(ram[3377]), .S(n12682), .Y(n8793) );
  MUX2X1 U10536 ( .B(ram[3329]), .A(ram[3345]), .S(n12645), .Y(n8792) );
  MUX2X1 U10537 ( .B(n8791), .A(n8788), .S(n12589), .Y(n8795) );
  MUX2X1 U10538 ( .B(ram[3297]), .A(ram[3313]), .S(n12640), .Y(n8799) );
  MUX2X1 U10539 ( .B(ram[3265]), .A(ram[3281]), .S(n12621), .Y(n8798) );
  MUX2X1 U10540 ( .B(ram[3233]), .A(ram[3249]), .S(n12664), .Y(n8802) );
  MUX2X1 U10541 ( .B(ram[3201]), .A(ram[3217]), .S(n12639), .Y(n8801) );
  MUX2X1 U10542 ( .B(n8800), .A(n8797), .S(n12586), .Y(n8811) );
  MUX2X1 U10543 ( .B(ram[3169]), .A(ram[3185]), .S(n12633), .Y(n8805) );
  MUX2X1 U10544 ( .B(ram[3137]), .A(ram[3153]), .S(n12643), .Y(n8804) );
  MUX2X1 U10545 ( .B(ram[3105]), .A(ram[3121]), .S(n12626), .Y(n8808) );
  MUX2X1 U10546 ( .B(ram[3073]), .A(ram[3089]), .S(n12640), .Y(n8807) );
  MUX2X1 U10547 ( .B(n8806), .A(n8803), .S(n12586), .Y(n8810) );
  MUX2X1 U10548 ( .B(n8809), .A(n8794), .S(n12566), .Y(n8813) );
  MUX2X1 U10549 ( .B(ram[3041]), .A(ram[3057]), .S(n12633), .Y(n8817) );
  MUX2X1 U10550 ( .B(ram[3009]), .A(ram[3025]), .S(n12645), .Y(n8816) );
  MUX2X1 U10551 ( .B(ram[2977]), .A(ram[2993]), .S(n12625), .Y(n8820) );
  MUX2X1 U10552 ( .B(ram[2945]), .A(ram[2961]), .S(n12629), .Y(n8819) );
  MUX2X1 U10553 ( .B(n8818), .A(n8815), .S(n12577), .Y(n8829) );
  MUX2X1 U10554 ( .B(ram[2913]), .A(ram[2929]), .S(n12651), .Y(n8823) );
  MUX2X1 U10555 ( .B(ram[2881]), .A(ram[2897]), .S(n12629), .Y(n8822) );
  MUX2X1 U10556 ( .B(ram[2849]), .A(ram[2865]), .S(n12629), .Y(n8826) );
  MUX2X1 U10557 ( .B(ram[2817]), .A(ram[2833]), .S(n12634), .Y(n8825) );
  MUX2X1 U10558 ( .B(n8824), .A(n8821), .S(n12582), .Y(n8828) );
  MUX2X1 U10559 ( .B(ram[2785]), .A(ram[2801]), .S(n12671), .Y(n8832) );
  MUX2X1 U10560 ( .B(ram[2753]), .A(ram[2769]), .S(n12638), .Y(n8831) );
  MUX2X1 U10561 ( .B(ram[2721]), .A(ram[2737]), .S(n12629), .Y(n8835) );
  MUX2X1 U10562 ( .B(ram[2689]), .A(ram[2705]), .S(n12638), .Y(n8834) );
  MUX2X1 U10563 ( .B(n8833), .A(n8830), .S(n12576), .Y(n8844) );
  MUX2X1 U10564 ( .B(ram[2657]), .A(ram[2673]), .S(n12674), .Y(n8838) );
  MUX2X1 U10565 ( .B(ram[2625]), .A(ram[2641]), .S(n12676), .Y(n8837) );
  MUX2X1 U10566 ( .B(ram[2593]), .A(ram[2609]), .S(n12671), .Y(n8841) );
  MUX2X1 U10567 ( .B(ram[2561]), .A(ram[2577]), .S(n12636), .Y(n8840) );
  MUX2X1 U10568 ( .B(n8839), .A(n8836), .S(n12579), .Y(n8843) );
  MUX2X1 U10569 ( .B(n8842), .A(n8827), .S(n12566), .Y(n8877) );
  MUX2X1 U10570 ( .B(ram[2529]), .A(ram[2545]), .S(n12652), .Y(n8847) );
  MUX2X1 U10571 ( .B(ram[2497]), .A(ram[2513]), .S(n12669), .Y(n8846) );
  MUX2X1 U10572 ( .B(ram[2465]), .A(ram[2481]), .S(n12631), .Y(n8850) );
  MUX2X1 U10573 ( .B(ram[2433]), .A(ram[2449]), .S(n12674), .Y(n8849) );
  MUX2X1 U10574 ( .B(n8848), .A(n8845), .S(n12586), .Y(n8859) );
  MUX2X1 U10575 ( .B(ram[2401]), .A(ram[2417]), .S(n12630), .Y(n8853) );
  MUX2X1 U10576 ( .B(ram[2369]), .A(ram[2385]), .S(n12672), .Y(n8852) );
  MUX2X1 U10577 ( .B(ram[2337]), .A(ram[2353]), .S(n12632), .Y(n8856) );
  MUX2X1 U10578 ( .B(ram[2305]), .A(ram[2321]), .S(n12661), .Y(n8855) );
  MUX2X1 U10579 ( .B(n8854), .A(n8851), .S(n12585), .Y(n8858) );
  MUX2X1 U10580 ( .B(ram[2273]), .A(ram[2289]), .S(n12632), .Y(n8862) );
  MUX2X1 U10581 ( .B(ram[2241]), .A(ram[2257]), .S(n12655), .Y(n8861) );
  MUX2X1 U10582 ( .B(ram[2209]), .A(ram[2225]), .S(n12633), .Y(n8865) );
  MUX2X1 U10583 ( .B(ram[2177]), .A(ram[2193]), .S(n12669), .Y(n8864) );
  MUX2X1 U10584 ( .B(n8863), .A(n8860), .S(n12587), .Y(n8874) );
  MUX2X1 U10585 ( .B(ram[2145]), .A(ram[2161]), .S(n12636), .Y(n8868) );
  MUX2X1 U10586 ( .B(ram[2113]), .A(ram[2129]), .S(n12680), .Y(n8867) );
  MUX2X1 U10587 ( .B(ram[2081]), .A(ram[2097]), .S(n12635), .Y(n8871) );
  MUX2X1 U10588 ( .B(ram[2049]), .A(ram[2065]), .S(n12621), .Y(n8870) );
  MUX2X1 U10589 ( .B(n8869), .A(n8866), .S(n12587), .Y(n8873) );
  MUX2X1 U10590 ( .B(n8872), .A(n8857), .S(n12565), .Y(n8876) );
  MUX2X1 U10591 ( .B(n8875), .A(n8812), .S(mem_access_addr[6]), .Y(n9005) );
  MUX2X1 U10592 ( .B(ram[2017]), .A(ram[2033]), .S(n12635), .Y(n8880) );
  MUX2X1 U10593 ( .B(ram[1985]), .A(ram[2001]), .S(n12667), .Y(n8879) );
  MUX2X1 U10594 ( .B(ram[1953]), .A(ram[1969]), .S(n12664), .Y(n8883) );
  MUX2X1 U10595 ( .B(ram[1921]), .A(ram[1937]), .S(n12650), .Y(n8882) );
  MUX2X1 U10596 ( .B(n8881), .A(n8878), .S(n12577), .Y(n8892) );
  MUX2X1 U10597 ( .B(ram[1889]), .A(ram[1905]), .S(n12678), .Y(n8886) );
  MUX2X1 U10598 ( .B(ram[1857]), .A(ram[1873]), .S(n12662), .Y(n8885) );
  MUX2X1 U10599 ( .B(ram[1825]), .A(ram[1841]), .S(n12683), .Y(n8889) );
  MUX2X1 U10600 ( .B(ram[1793]), .A(ram[1809]), .S(n12625), .Y(n8888) );
  MUX2X1 U10601 ( .B(n8887), .A(n8884), .S(n12589), .Y(n8891) );
  MUX2X1 U10602 ( .B(ram[1761]), .A(ram[1777]), .S(n12632), .Y(n8895) );
  MUX2X1 U10603 ( .B(ram[1729]), .A(ram[1745]), .S(n12666), .Y(n8894) );
  MUX2X1 U10604 ( .B(ram[1697]), .A(ram[1713]), .S(n12631), .Y(n8898) );
  MUX2X1 U10605 ( .B(ram[1665]), .A(ram[1681]), .S(n12658), .Y(n8897) );
  MUX2X1 U10606 ( .B(n8896), .A(n8893), .S(n12581), .Y(n8907) );
  MUX2X1 U10607 ( .B(ram[1633]), .A(ram[1649]), .S(n12626), .Y(n8901) );
  MUX2X1 U10608 ( .B(ram[1601]), .A(ram[1617]), .S(n12681), .Y(n8900) );
  MUX2X1 U10609 ( .B(ram[1569]), .A(ram[1585]), .S(mem_access_addr[0]), .Y(
        n8904) );
  MUX2X1 U10610 ( .B(ram[1537]), .A(ram[1553]), .S(n12649), .Y(n8903) );
  MUX2X1 U10611 ( .B(n8902), .A(n8899), .S(n12586), .Y(n8906) );
  MUX2X1 U10612 ( .B(n8905), .A(n8890), .S(n12566), .Y(n8940) );
  MUX2X1 U10613 ( .B(ram[1505]), .A(ram[1521]), .S(n12648), .Y(n8910) );
  MUX2X1 U10614 ( .B(ram[1473]), .A(ram[1489]), .S(n12662), .Y(n8909) );
  MUX2X1 U10615 ( .B(ram[1441]), .A(ram[1457]), .S(n12682), .Y(n8913) );
  MUX2X1 U10616 ( .B(ram[1409]), .A(ram[1425]), .S(n12651), .Y(n8912) );
  MUX2X1 U10617 ( .B(n8911), .A(n8908), .S(n12582), .Y(n8922) );
  MUX2X1 U10618 ( .B(ram[1377]), .A(ram[1393]), .S(n12668), .Y(n8916) );
  MUX2X1 U10619 ( .B(ram[1345]), .A(ram[1361]), .S(n12640), .Y(n8915) );
  MUX2X1 U10620 ( .B(ram[1313]), .A(ram[1329]), .S(n12676), .Y(n8919) );
  MUX2X1 U10621 ( .B(ram[1281]), .A(ram[1297]), .S(n12667), .Y(n8918) );
  MUX2X1 U10622 ( .B(n8917), .A(n8914), .S(n12589), .Y(n8921) );
  MUX2X1 U10623 ( .B(ram[1249]), .A(ram[1265]), .S(n12656), .Y(n8925) );
  MUX2X1 U10624 ( .B(ram[1217]), .A(ram[1233]), .S(n12625), .Y(n8924) );
  MUX2X1 U10625 ( .B(ram[1185]), .A(ram[1201]), .S(n12671), .Y(n8928) );
  MUX2X1 U10626 ( .B(ram[1153]), .A(ram[1169]), .S(n12676), .Y(n8927) );
  MUX2X1 U10627 ( .B(n8926), .A(n8923), .S(mem_access_addr[2]), .Y(n8937) );
  MUX2X1 U10628 ( .B(ram[1121]), .A(ram[1137]), .S(n12683), .Y(n8931) );
  MUX2X1 U10629 ( .B(ram[1089]), .A(ram[1105]), .S(n12624), .Y(n8930) );
  MUX2X1 U10630 ( .B(ram[1057]), .A(ram[1073]), .S(n12663), .Y(n8934) );
  MUX2X1 U10631 ( .B(ram[1025]), .A(ram[1041]), .S(n12648), .Y(n8933) );
  MUX2X1 U10632 ( .B(n8932), .A(n8929), .S(n12583), .Y(n8936) );
  MUX2X1 U10633 ( .B(n8935), .A(n8920), .S(n12565), .Y(n8939) );
  MUX2X1 U10634 ( .B(ram[993]), .A(ram[1009]), .S(n12668), .Y(n8943) );
  MUX2X1 U10635 ( .B(ram[961]), .A(ram[977]), .S(n12653), .Y(n8942) );
  MUX2X1 U10636 ( .B(ram[929]), .A(ram[945]), .S(n12627), .Y(n8946) );
  MUX2X1 U10637 ( .B(ram[897]), .A(ram[913]), .S(n12642), .Y(n8945) );
  MUX2X1 U10638 ( .B(n8944), .A(n8941), .S(n12579), .Y(n8955) );
  MUX2X1 U10639 ( .B(ram[865]), .A(ram[881]), .S(n12664), .Y(n8949) );
  MUX2X1 U10640 ( .B(ram[833]), .A(ram[849]), .S(n12624), .Y(n8948) );
  MUX2X1 U10641 ( .B(ram[801]), .A(ram[817]), .S(n12642), .Y(n8952) );
  MUX2X1 U10642 ( .B(ram[769]), .A(ram[785]), .S(n12669), .Y(n8951) );
  MUX2X1 U10643 ( .B(n8950), .A(n8947), .S(n12578), .Y(n8954) );
  MUX2X1 U10644 ( .B(ram[737]), .A(ram[753]), .S(n12673), .Y(n8958) );
  MUX2X1 U10645 ( .B(ram[705]), .A(ram[721]), .S(n12623), .Y(n8957) );
  MUX2X1 U10646 ( .B(ram[673]), .A(ram[689]), .S(n12629), .Y(n8961) );
  MUX2X1 U10647 ( .B(ram[641]), .A(ram[657]), .S(n12652), .Y(n8960) );
  MUX2X1 U10648 ( .B(n8959), .A(n8956), .S(n12583), .Y(n8970) );
  MUX2X1 U10649 ( .B(ram[609]), .A(ram[625]), .S(n12661), .Y(n8964) );
  MUX2X1 U10650 ( .B(ram[577]), .A(ram[593]), .S(n12641), .Y(n8963) );
  MUX2X1 U10651 ( .B(ram[545]), .A(ram[561]), .S(n12671), .Y(n8967) );
  MUX2X1 U10652 ( .B(ram[513]), .A(ram[529]), .S(n12624), .Y(n8966) );
  MUX2X1 U10653 ( .B(n8965), .A(n8962), .S(n12583), .Y(n8969) );
  MUX2X1 U10654 ( .B(n8968), .A(n8953), .S(n12565), .Y(n9003) );
  MUX2X1 U10655 ( .B(ram[481]), .A(ram[497]), .S(n12672), .Y(n8973) );
  MUX2X1 U10656 ( .B(ram[449]), .A(ram[465]), .S(n12654), .Y(n8972) );
  MUX2X1 U10657 ( .B(ram[417]), .A(ram[433]), .S(n12668), .Y(n8976) );
  MUX2X1 U10658 ( .B(ram[385]), .A(ram[401]), .S(n12682), .Y(n8975) );
  MUX2X1 U10659 ( .B(n8974), .A(n8971), .S(n12588), .Y(n8985) );
  MUX2X1 U10660 ( .B(ram[353]), .A(ram[369]), .S(mem_access_addr[0]), .Y(n8979) );
  MUX2X1 U10661 ( .B(ram[321]), .A(ram[337]), .S(n12670), .Y(n8978) );
  MUX2X1 U10662 ( .B(ram[289]), .A(ram[305]), .S(n12669), .Y(n8982) );
  MUX2X1 U10663 ( .B(ram[257]), .A(ram[273]), .S(n12683), .Y(n8981) );
  MUX2X1 U10664 ( .B(n8980), .A(n8977), .S(n12577), .Y(n8984) );
  MUX2X1 U10665 ( .B(ram[225]), .A(ram[241]), .S(n12623), .Y(n8988) );
  MUX2X1 U10666 ( .B(ram[193]), .A(ram[209]), .S(n12667), .Y(n8987) );
  MUX2X1 U10667 ( .B(ram[161]), .A(ram[177]), .S(n12628), .Y(n8991) );
  MUX2X1 U10668 ( .B(ram[129]), .A(ram[145]), .S(n12634), .Y(n8990) );
  MUX2X1 U10669 ( .B(n8989), .A(n8986), .S(n12579), .Y(n9000) );
  MUX2X1 U10670 ( .B(ram[97]), .A(ram[113]), .S(n12679), .Y(n8994) );
  MUX2X1 U10671 ( .B(ram[65]), .A(ram[81]), .S(n12683), .Y(n8993) );
  MUX2X1 U10672 ( .B(ram[33]), .A(ram[49]), .S(mem_access_addr[0]), .Y(n8997)
         );
  MUX2X1 U10673 ( .B(ram[1]), .A(ram[17]), .S(n12677), .Y(n8996) );
  MUX2X1 U10674 ( .B(n8995), .A(n8992), .S(n12578), .Y(n8999) );
  MUX2X1 U10675 ( .B(n8998), .A(n8983), .S(n12566), .Y(n9002) );
  MUX2X1 U10676 ( .B(n9001), .A(n8938), .S(n1), .Y(n9004) );
  MUX2X1 U10677 ( .B(ram[4066]), .A(ram[4082]), .S(n12622), .Y(n9008) );
  MUX2X1 U10678 ( .B(ram[4034]), .A(ram[4050]), .S(n12683), .Y(n9007) );
  MUX2X1 U10679 ( .B(ram[4002]), .A(ram[4018]), .S(n12624), .Y(n9011) );
  MUX2X1 U10680 ( .B(ram[3970]), .A(ram[3986]), .S(n12683), .Y(n9010) );
  MUX2X1 U10681 ( .B(n9009), .A(n9006), .S(n12577), .Y(n9020) );
  MUX2X1 U10682 ( .B(ram[3938]), .A(ram[3954]), .S(n12631), .Y(n9014) );
  MUX2X1 U10683 ( .B(ram[3906]), .A(ram[3922]), .S(n12683), .Y(n9013) );
  MUX2X1 U10684 ( .B(ram[3874]), .A(ram[3890]), .S(n12678), .Y(n9017) );
  MUX2X1 U10685 ( .B(ram[3842]), .A(ram[3858]), .S(n12654), .Y(n9016) );
  MUX2X1 U10686 ( .B(n9015), .A(n9012), .S(n12584), .Y(n9019) );
  MUX2X1 U10687 ( .B(ram[3810]), .A(ram[3826]), .S(n12632), .Y(n9023) );
  MUX2X1 U10688 ( .B(ram[3778]), .A(ram[3794]), .S(n12634), .Y(n9022) );
  MUX2X1 U10689 ( .B(ram[3746]), .A(ram[3762]), .S(n12626), .Y(n9026) );
  MUX2X1 U10690 ( .B(ram[3714]), .A(ram[3730]), .S(n12629), .Y(n9025) );
  MUX2X1 U10691 ( .B(n9024), .A(n9021), .S(n12575), .Y(n9035) );
  MUX2X1 U10692 ( .B(ram[3682]), .A(ram[3698]), .S(n12628), .Y(n9029) );
  MUX2X1 U10693 ( .B(ram[3650]), .A(ram[3666]), .S(n12669), .Y(n9028) );
  MUX2X1 U10694 ( .B(ram[3618]), .A(ram[3634]), .S(n12654), .Y(n9032) );
  MUX2X1 U10695 ( .B(ram[3586]), .A(ram[3602]), .S(n12641), .Y(n9031) );
  MUX2X1 U10696 ( .B(n9030), .A(n9027), .S(n12575), .Y(n9034) );
  MUX2X1 U10697 ( .B(n9033), .A(n9018), .S(n12566), .Y(n9068) );
  MUX2X1 U10698 ( .B(ram[3554]), .A(ram[3570]), .S(n12622), .Y(n9038) );
  MUX2X1 U10699 ( .B(ram[3522]), .A(ram[3538]), .S(n12635), .Y(n9037) );
  MUX2X1 U10700 ( .B(ram[3490]), .A(ram[3506]), .S(n12677), .Y(n9041) );
  MUX2X1 U10701 ( .B(ram[3458]), .A(ram[3474]), .S(n12623), .Y(n9040) );
  MUX2X1 U10702 ( .B(n9039), .A(n9036), .S(n12588), .Y(n9050) );
  MUX2X1 U10703 ( .B(ram[3426]), .A(ram[3442]), .S(n12670), .Y(n9044) );
  MUX2X1 U10704 ( .B(ram[3394]), .A(ram[3410]), .S(n12654), .Y(n9043) );
  MUX2X1 U10705 ( .B(ram[3362]), .A(ram[3378]), .S(n12646), .Y(n9047) );
  MUX2X1 U10706 ( .B(ram[3330]), .A(ram[3346]), .S(n12629), .Y(n9046) );
  MUX2X1 U10707 ( .B(n9045), .A(n9042), .S(n12579), .Y(n9049) );
  MUX2X1 U10708 ( .B(ram[3298]), .A(ram[3314]), .S(n12679), .Y(n9053) );
  MUX2X1 U10709 ( .B(ram[3266]), .A(ram[3282]), .S(n12663), .Y(n9052) );
  MUX2X1 U10710 ( .B(ram[3234]), .A(ram[3250]), .S(n12639), .Y(n9056) );
  MUX2X1 U10711 ( .B(ram[3202]), .A(ram[3218]), .S(n12680), .Y(n9055) );
  MUX2X1 U10712 ( .B(n9054), .A(n9051), .S(n12579), .Y(n9065) );
  MUX2X1 U10713 ( .B(ram[3170]), .A(ram[3186]), .S(n12658), .Y(n9059) );
  MUX2X1 U10714 ( .B(ram[3138]), .A(ram[3154]), .S(n12676), .Y(n9058) );
  MUX2X1 U10715 ( .B(ram[3106]), .A(ram[3122]), .S(n12624), .Y(n9062) );
  MUX2X1 U10716 ( .B(ram[3074]), .A(ram[3090]), .S(n12674), .Y(n9061) );
  MUX2X1 U10717 ( .B(n9060), .A(n9057), .S(n12582), .Y(n9064) );
  MUX2X1 U10718 ( .B(n9063), .A(n9048), .S(n12565), .Y(n9067) );
  MUX2X1 U10719 ( .B(ram[3042]), .A(ram[3058]), .S(n12639), .Y(n9071) );
  MUX2X1 U10720 ( .B(ram[3010]), .A(ram[3026]), .S(n12662), .Y(n9070) );
  MUX2X1 U10721 ( .B(ram[2978]), .A(ram[2994]), .S(n12639), .Y(n9074) );
  MUX2X1 U10722 ( .B(ram[2946]), .A(ram[2962]), .S(n12632), .Y(n9073) );
  MUX2X1 U10723 ( .B(n9072), .A(n9069), .S(n12588), .Y(n9083) );
  MUX2X1 U10724 ( .B(ram[2914]), .A(ram[2930]), .S(n12682), .Y(n9077) );
  MUX2X1 U10725 ( .B(ram[2882]), .A(ram[2898]), .S(mem_access_addr[0]), .Y(
        n9076) );
  MUX2X1 U10726 ( .B(ram[2850]), .A(ram[2866]), .S(n12680), .Y(n9080) );
  MUX2X1 U10727 ( .B(ram[2818]), .A(ram[2834]), .S(n12679), .Y(n9079) );
  MUX2X1 U10728 ( .B(n9078), .A(n9075), .S(n12589), .Y(n9082) );
  MUX2X1 U10729 ( .B(ram[2786]), .A(ram[2802]), .S(n12630), .Y(n9086) );
  MUX2X1 U10730 ( .B(ram[2754]), .A(ram[2770]), .S(n12682), .Y(n9085) );
  MUX2X1 U10731 ( .B(ram[2722]), .A(ram[2738]), .S(n12666), .Y(n9089) );
  MUX2X1 U10732 ( .B(ram[2690]), .A(ram[2706]), .S(n12632), .Y(n9088) );
  MUX2X1 U10733 ( .B(n9087), .A(n9084), .S(n12587), .Y(n9098) );
  MUX2X1 U10734 ( .B(ram[2658]), .A(ram[2674]), .S(n12630), .Y(n9092) );
  MUX2X1 U10735 ( .B(ram[2626]), .A(ram[2642]), .S(n12654), .Y(n9091) );
  MUX2X1 U10736 ( .B(ram[2594]), .A(ram[2610]), .S(n12633), .Y(n9095) );
  MUX2X1 U10737 ( .B(ram[2562]), .A(ram[2578]), .S(n12664), .Y(n9094) );
  MUX2X1 U10738 ( .B(n9093), .A(n9090), .S(n12582), .Y(n9097) );
  MUX2X1 U10739 ( .B(n9096), .A(n9081), .S(n12567), .Y(n9131) );
  MUX2X1 U10740 ( .B(ram[2530]), .A(ram[2546]), .S(n12681), .Y(n9101) );
  MUX2X1 U10741 ( .B(ram[2498]), .A(ram[2514]), .S(n12673), .Y(n9100) );
  MUX2X1 U10742 ( .B(ram[2466]), .A(ram[2482]), .S(n12630), .Y(n9104) );
  MUX2X1 U10743 ( .B(ram[2434]), .A(ram[2450]), .S(n12665), .Y(n9103) );
  MUX2X1 U10744 ( .B(n9102), .A(n9099), .S(n12589), .Y(n9113) );
  MUX2X1 U10745 ( .B(ram[2402]), .A(ram[2418]), .S(n12622), .Y(n9107) );
  MUX2X1 U10746 ( .B(ram[2370]), .A(ram[2386]), .S(n12676), .Y(n9106) );
  MUX2X1 U10747 ( .B(ram[2338]), .A(ram[2354]), .S(n12658), .Y(n9110) );
  MUX2X1 U10748 ( .B(ram[2306]), .A(ram[2322]), .S(n12667), .Y(n9109) );
  MUX2X1 U10749 ( .B(n9108), .A(n9105), .S(n12581), .Y(n9112) );
  MUX2X1 U10750 ( .B(ram[2274]), .A(ram[2290]), .S(n12664), .Y(n9116) );
  MUX2X1 U10751 ( .B(ram[2242]), .A(ram[2258]), .S(n12622), .Y(n9115) );
  MUX2X1 U10752 ( .B(ram[2210]), .A(ram[2226]), .S(n12653), .Y(n9119) );
  MUX2X1 U10753 ( .B(ram[2178]), .A(ram[2194]), .S(n12630), .Y(n9118) );
  MUX2X1 U10754 ( .B(n9117), .A(n9114), .S(n12586), .Y(n9128) );
  MUX2X1 U10755 ( .B(ram[2146]), .A(ram[2162]), .S(n12624), .Y(n9122) );
  MUX2X1 U10756 ( .B(ram[2114]), .A(ram[2130]), .S(mem_access_addr[0]), .Y(
        n9121) );
  MUX2X1 U10757 ( .B(ram[2082]), .A(ram[2098]), .S(n12627), .Y(n9125) );
  MUX2X1 U10758 ( .B(ram[2050]), .A(ram[2066]), .S(n12662), .Y(n9124) );
  MUX2X1 U10759 ( .B(n9123), .A(n9120), .S(n12576), .Y(n9127) );
  MUX2X1 U10760 ( .B(n9126), .A(n9111), .S(n12567), .Y(n9130) );
  MUX2X1 U10761 ( .B(n9129), .A(n9066), .S(mem_access_addr[6]), .Y(n9259) );
  MUX2X1 U10762 ( .B(ram[2018]), .A(ram[2034]), .S(n12678), .Y(n9134) );
  MUX2X1 U10763 ( .B(ram[1986]), .A(ram[2002]), .S(n12636), .Y(n9133) );
  MUX2X1 U10764 ( .B(ram[1954]), .A(ram[1970]), .S(n12680), .Y(n9137) );
  MUX2X1 U10765 ( .B(ram[1922]), .A(ram[1938]), .S(n12633), .Y(n9136) );
  MUX2X1 U10766 ( .B(n9135), .A(n9132), .S(n12577), .Y(n9146) );
  MUX2X1 U10767 ( .B(ram[1890]), .A(ram[1906]), .S(n12639), .Y(n9140) );
  MUX2X1 U10768 ( .B(ram[1858]), .A(ram[1874]), .S(n12634), .Y(n9139) );
  MUX2X1 U10769 ( .B(ram[1826]), .A(ram[1842]), .S(n12621), .Y(n9143) );
  MUX2X1 U10770 ( .B(ram[1794]), .A(ram[1810]), .S(n12642), .Y(n9142) );
  MUX2X1 U10771 ( .B(n9141), .A(n9138), .S(n12589), .Y(n9145) );
  MUX2X1 U10772 ( .B(ram[1762]), .A(ram[1778]), .S(n12663), .Y(n9149) );
  MUX2X1 U10773 ( .B(ram[1730]), .A(ram[1746]), .S(n12668), .Y(n9148) );
  MUX2X1 U10774 ( .B(ram[1698]), .A(ram[1714]), .S(n12653), .Y(n9152) );
  MUX2X1 U10775 ( .B(ram[1666]), .A(ram[1682]), .S(n12655), .Y(n9151) );
  MUX2X1 U10776 ( .B(n9150), .A(n9147), .S(n12575), .Y(n9161) );
  MUX2X1 U10777 ( .B(ram[1634]), .A(ram[1650]), .S(n12622), .Y(n9155) );
  MUX2X1 U10778 ( .B(ram[1602]), .A(ram[1618]), .S(n12651), .Y(n9154) );
  MUX2X1 U10779 ( .B(ram[1570]), .A(ram[1586]), .S(n12682), .Y(n9158) );
  MUX2X1 U10780 ( .B(ram[1538]), .A(ram[1554]), .S(n12641), .Y(n9157) );
  MUX2X1 U10781 ( .B(n9156), .A(n9153), .S(mem_access_addr[2]), .Y(n9160) );
  MUX2X1 U10782 ( .B(n9159), .A(n9144), .S(n12567), .Y(n9194) );
  MUX2X1 U10783 ( .B(ram[1506]), .A(ram[1522]), .S(mem_access_addr[0]), .Y(
        n9164) );
  MUX2X1 U10784 ( .B(ram[1474]), .A(ram[1490]), .S(n12644), .Y(n9163) );
  MUX2X1 U10785 ( .B(ram[1442]), .A(ram[1458]), .S(n12652), .Y(n9167) );
  MUX2X1 U10786 ( .B(ram[1410]), .A(ram[1426]), .S(n12643), .Y(n9166) );
  MUX2X1 U10787 ( .B(n9165), .A(n9162), .S(n12589), .Y(n9176) );
  MUX2X1 U10788 ( .B(ram[1378]), .A(ram[1394]), .S(n12639), .Y(n9170) );
  MUX2X1 U10789 ( .B(ram[1346]), .A(ram[1362]), .S(n12682), .Y(n9169) );
  MUX2X1 U10790 ( .B(ram[1314]), .A(ram[1330]), .S(n12644), .Y(n9173) );
  MUX2X1 U10791 ( .B(ram[1282]), .A(ram[1298]), .S(n12640), .Y(n9172) );
  MUX2X1 U10792 ( .B(n9171), .A(n9168), .S(n12579), .Y(n9175) );
  MUX2X1 U10793 ( .B(ram[1250]), .A(ram[1266]), .S(n12650), .Y(n9179) );
  MUX2X1 U10794 ( .B(ram[1218]), .A(ram[1234]), .S(n12663), .Y(n9178) );
  MUX2X1 U10795 ( .B(ram[1186]), .A(ram[1202]), .S(n12637), .Y(n9182) );
  MUX2X1 U10796 ( .B(ram[1154]), .A(ram[1170]), .S(n12663), .Y(n9181) );
  MUX2X1 U10797 ( .B(n9180), .A(n9177), .S(n12578), .Y(n9191) );
  MUX2X1 U10798 ( .B(ram[1122]), .A(ram[1138]), .S(n12683), .Y(n9185) );
  MUX2X1 U10799 ( .B(ram[1090]), .A(ram[1106]), .S(n12626), .Y(n9184) );
  MUX2X1 U10800 ( .B(ram[1058]), .A(ram[1074]), .S(n12672), .Y(n9188) );
  MUX2X1 U10801 ( .B(ram[1026]), .A(ram[1042]), .S(n12628), .Y(n9187) );
  MUX2X1 U10802 ( .B(n9186), .A(n9183), .S(n12578), .Y(n9190) );
  MUX2X1 U10803 ( .B(n9189), .A(n9174), .S(n12567), .Y(n9193) );
  MUX2X1 U10804 ( .B(ram[994]), .A(ram[1010]), .S(n12621), .Y(n9197) );
  MUX2X1 U10805 ( .B(ram[962]), .A(ram[978]), .S(n12661), .Y(n9196) );
  MUX2X1 U10806 ( .B(ram[930]), .A(ram[946]), .S(n12632), .Y(n9200) );
  MUX2X1 U10807 ( .B(ram[898]), .A(ram[914]), .S(n12622), .Y(n9199) );
  MUX2X1 U10808 ( .B(n9198), .A(n9195), .S(n12577), .Y(n9209) );
  MUX2X1 U10809 ( .B(ram[866]), .A(ram[882]), .S(n12633), .Y(n9203) );
  MUX2X1 U10810 ( .B(ram[834]), .A(ram[850]), .S(n12669), .Y(n9202) );
  MUX2X1 U10811 ( .B(ram[802]), .A(ram[818]), .S(n12631), .Y(n9206) );
  MUX2X1 U10812 ( .B(ram[770]), .A(ram[786]), .S(n12647), .Y(n9205) );
  MUX2X1 U10813 ( .B(n9204), .A(n9201), .S(n12588), .Y(n9208) );
  MUX2X1 U10814 ( .B(ram[738]), .A(ram[754]), .S(n12625), .Y(n9212) );
  MUX2X1 U10815 ( .B(ram[706]), .A(ram[722]), .S(n12629), .Y(n9211) );
  MUX2X1 U10816 ( .B(ram[674]), .A(ram[690]), .S(n12636), .Y(n9215) );
  MUX2X1 U10817 ( .B(ram[642]), .A(ram[658]), .S(n12633), .Y(n9214) );
  MUX2X1 U10818 ( .B(n9213), .A(n9210), .S(n12575), .Y(n9224) );
  MUX2X1 U10819 ( .B(ram[610]), .A(ram[626]), .S(n12681), .Y(n9218) );
  MUX2X1 U10820 ( .B(ram[578]), .A(ram[594]), .S(n12656), .Y(n9217) );
  MUX2X1 U10821 ( .B(ram[546]), .A(ram[562]), .S(n12632), .Y(n9221) );
  MUX2X1 U10822 ( .B(ram[514]), .A(ram[530]), .S(n12646), .Y(n9220) );
  MUX2X1 U10823 ( .B(n9219), .A(n9216), .S(n12575), .Y(n9223) );
  MUX2X1 U10824 ( .B(n9222), .A(n9207), .S(n12567), .Y(n9257) );
  MUX2X1 U10825 ( .B(ram[482]), .A(ram[498]), .S(n12621), .Y(n9227) );
  MUX2X1 U10826 ( .B(ram[450]), .A(ram[466]), .S(n12626), .Y(n9226) );
  MUX2X1 U10827 ( .B(ram[418]), .A(ram[434]), .S(n12639), .Y(n9230) );
  MUX2X1 U10828 ( .B(ram[386]), .A(ram[402]), .S(n12651), .Y(n9229) );
  MUX2X1 U10829 ( .B(n9228), .A(n9225), .S(n12586), .Y(n9239) );
  MUX2X1 U10830 ( .B(ram[354]), .A(ram[370]), .S(n12641), .Y(n9233) );
  MUX2X1 U10831 ( .B(ram[322]), .A(ram[338]), .S(n12662), .Y(n9232) );
  MUX2X1 U10832 ( .B(ram[290]), .A(ram[306]), .S(mem_access_addr[0]), .Y(n9236) );
  MUX2X1 U10833 ( .B(ram[258]), .A(ram[274]), .S(n12651), .Y(n9235) );
  MUX2X1 U10834 ( .B(n9234), .A(n9231), .S(n12588), .Y(n9238) );
  MUX2X1 U10835 ( .B(ram[226]), .A(ram[242]), .S(n12631), .Y(n9242) );
  MUX2X1 U10836 ( .B(ram[194]), .A(ram[210]), .S(n12656), .Y(n9241) );
  MUX2X1 U10837 ( .B(ram[162]), .A(ram[178]), .S(n12656), .Y(n9245) );
  MUX2X1 U10838 ( .B(ram[130]), .A(ram[146]), .S(n12682), .Y(n9244) );
  MUX2X1 U10839 ( .B(n9243), .A(n9240), .S(n12588), .Y(n9254) );
  MUX2X1 U10840 ( .B(ram[98]), .A(ram[114]), .S(n12641), .Y(n9248) );
  MUX2X1 U10841 ( .B(ram[66]), .A(ram[82]), .S(n12631), .Y(n9247) );
  MUX2X1 U10842 ( .B(ram[34]), .A(ram[50]), .S(n12667), .Y(n9251) );
  MUX2X1 U10843 ( .B(ram[2]), .A(ram[18]), .S(n12670), .Y(n9250) );
  MUX2X1 U10844 ( .B(n9249), .A(n9246), .S(n12589), .Y(n9253) );
  MUX2X1 U10845 ( .B(n9252), .A(n9237), .S(n12564), .Y(n9256) );
  MUX2X1 U10846 ( .B(n9255), .A(n9192), .S(mem_access_addr[6]), .Y(n9258) );
  MUX2X1 U10847 ( .B(ram[4067]), .A(ram[4083]), .S(n12674), .Y(n9262) );
  MUX2X1 U10848 ( .B(ram[4035]), .A(ram[4051]), .S(n12658), .Y(n9261) );
  MUX2X1 U10849 ( .B(ram[4003]), .A(ram[4019]), .S(n12637), .Y(n9265) );
  MUX2X1 U10850 ( .B(ram[3971]), .A(ram[3987]), .S(n12636), .Y(n9264) );
  MUX2X1 U10851 ( .B(n9263), .A(n9260), .S(n12581), .Y(n9274) );
  MUX2X1 U10852 ( .B(ram[3939]), .A(ram[3955]), .S(n12674), .Y(n9268) );
  MUX2X1 U10853 ( .B(ram[3907]), .A(ram[3923]), .S(n12671), .Y(n9267) );
  MUX2X1 U10854 ( .B(ram[3875]), .A(ram[3891]), .S(n12634), .Y(n9271) );
  MUX2X1 U10855 ( .B(ram[3843]), .A(ram[3859]), .S(n12681), .Y(n9270) );
  MUX2X1 U10856 ( .B(n9269), .A(n9266), .S(n12582), .Y(n9273) );
  MUX2X1 U10857 ( .B(ram[3811]), .A(ram[3827]), .S(n12633), .Y(n9277) );
  MUX2X1 U10858 ( .B(ram[3779]), .A(ram[3795]), .S(n12682), .Y(n9276) );
  MUX2X1 U10859 ( .B(ram[3747]), .A(ram[3763]), .S(n12682), .Y(n9280) );
  MUX2X1 U10860 ( .B(ram[3715]), .A(ram[3731]), .S(n12627), .Y(n9279) );
  MUX2X1 U10861 ( .B(n9278), .A(n9275), .S(n12589), .Y(n9289) );
  MUX2X1 U10862 ( .B(ram[3683]), .A(ram[3699]), .S(n12664), .Y(n9283) );
  MUX2X1 U10863 ( .B(ram[3651]), .A(ram[3667]), .S(n12647), .Y(n9282) );
  MUX2X1 U10864 ( .B(ram[3619]), .A(ram[3635]), .S(n12663), .Y(n9286) );
  MUX2X1 U10865 ( .B(ram[3587]), .A(ram[3603]), .S(n12666), .Y(n9285) );
  MUX2X1 U10866 ( .B(n9284), .A(n9281), .S(n12580), .Y(n9288) );
  MUX2X1 U10867 ( .B(n9287), .A(n9272), .S(n12565), .Y(n9322) );
  MUX2X1 U10868 ( .B(ram[3555]), .A(ram[3571]), .S(n12654), .Y(n9292) );
  MUX2X1 U10869 ( .B(ram[3523]), .A(ram[3539]), .S(n12636), .Y(n9291) );
  MUX2X1 U10870 ( .B(ram[3491]), .A(ram[3507]), .S(n12664), .Y(n9295) );
  MUX2X1 U10871 ( .B(ram[3459]), .A(ram[3475]), .S(n12655), .Y(n9294) );
  MUX2X1 U10872 ( .B(n9293), .A(n9290), .S(n12586), .Y(n9304) );
  MUX2X1 U10873 ( .B(ram[3427]), .A(ram[3443]), .S(n12630), .Y(n9298) );
  MUX2X1 U10874 ( .B(ram[3395]), .A(ram[3411]), .S(n12621), .Y(n9297) );
  MUX2X1 U10875 ( .B(ram[3363]), .A(ram[3379]), .S(n12649), .Y(n9301) );
  MUX2X1 U10876 ( .B(ram[3331]), .A(ram[3347]), .S(n12647), .Y(n9300) );
  MUX2X1 U10877 ( .B(n9299), .A(n9296), .S(n12583), .Y(n9303) );
  MUX2X1 U10878 ( .B(ram[3299]), .A(ram[3315]), .S(n12667), .Y(n9307) );
  MUX2X1 U10879 ( .B(ram[3267]), .A(ram[3283]), .S(n12641), .Y(n9306) );
  MUX2X1 U10880 ( .B(ram[3235]), .A(ram[3251]), .S(n12632), .Y(n9310) );
  MUX2X1 U10881 ( .B(ram[3203]), .A(ram[3219]), .S(n12658), .Y(n9309) );
  MUX2X1 U10882 ( .B(n9308), .A(n9305), .S(n12586), .Y(n9319) );
  MUX2X1 U10883 ( .B(ram[3171]), .A(ram[3187]), .S(n12675), .Y(n9313) );
  MUX2X1 U10884 ( .B(ram[3139]), .A(ram[3155]), .S(n12661), .Y(n9312) );
  MUX2X1 U10885 ( .B(ram[3107]), .A(ram[3123]), .S(n12659), .Y(n9316) );
  MUX2X1 U10886 ( .B(ram[3075]), .A(ram[3091]), .S(n12670), .Y(n9315) );
  MUX2X1 U10887 ( .B(n9314), .A(n9311), .S(n12575), .Y(n9318) );
  MUX2X1 U10888 ( .B(n9317), .A(n9302), .S(n12564), .Y(n9321) );
  MUX2X1 U10889 ( .B(ram[3043]), .A(ram[3059]), .S(n12638), .Y(n9325) );
  MUX2X1 U10890 ( .B(ram[3011]), .A(ram[3027]), .S(n12683), .Y(n9324) );
  MUX2X1 U10891 ( .B(ram[2979]), .A(ram[2995]), .S(n12625), .Y(n9328) );
  MUX2X1 U10892 ( .B(ram[2947]), .A(ram[2963]), .S(n12628), .Y(n9327) );
  MUX2X1 U10893 ( .B(n9326), .A(n9323), .S(n12587), .Y(n9337) );
  MUX2X1 U10894 ( .B(ram[2915]), .A(ram[2931]), .S(n12628), .Y(n9331) );
  MUX2X1 U10895 ( .B(ram[2883]), .A(ram[2899]), .S(n12678), .Y(n9330) );
  MUX2X1 U10896 ( .B(ram[2851]), .A(ram[2867]), .S(n12653), .Y(n9334) );
  MUX2X1 U10897 ( .B(ram[2819]), .A(ram[2835]), .S(n12635), .Y(n9333) );
  MUX2X1 U10898 ( .B(n9332), .A(n9329), .S(n12588), .Y(n9336) );
  MUX2X1 U10899 ( .B(ram[2787]), .A(ram[2803]), .S(n12635), .Y(n9340) );
  MUX2X1 U10900 ( .B(ram[2755]), .A(ram[2771]), .S(n12637), .Y(n9339) );
  MUX2X1 U10901 ( .B(ram[2723]), .A(ram[2739]), .S(n12635), .Y(n9343) );
  MUX2X1 U10902 ( .B(ram[2691]), .A(ram[2707]), .S(n12649), .Y(n9342) );
  MUX2X1 U10903 ( .B(n9341), .A(n9338), .S(n12589), .Y(n9352) );
  MUX2X1 U10904 ( .B(ram[2659]), .A(ram[2675]), .S(n12633), .Y(n9346) );
  MUX2X1 U10905 ( .B(ram[2627]), .A(ram[2643]), .S(n12627), .Y(n9345) );
  MUX2X1 U10906 ( .B(ram[2595]), .A(ram[2611]), .S(n12625), .Y(n9349) );
  MUX2X1 U10907 ( .B(ram[2563]), .A(ram[2579]), .S(n12678), .Y(n9348) );
  MUX2X1 U10908 ( .B(n9347), .A(n9344), .S(n12587), .Y(n9351) );
  MUX2X1 U10909 ( .B(n9350), .A(n9335), .S(n12564), .Y(n9385) );
  MUX2X1 U10910 ( .B(ram[2531]), .A(ram[2547]), .S(n12650), .Y(n9355) );
  MUX2X1 U10911 ( .B(ram[2499]), .A(ram[2515]), .S(n12621), .Y(n9354) );
  MUX2X1 U10912 ( .B(ram[2467]), .A(ram[2483]), .S(n12642), .Y(n9358) );
  MUX2X1 U10913 ( .B(ram[2435]), .A(ram[2451]), .S(n12661), .Y(n9357) );
  MUX2X1 U10914 ( .B(n9356), .A(n9353), .S(n12588), .Y(n9367) );
  MUX2X1 U10915 ( .B(ram[2403]), .A(ram[2419]), .S(n12643), .Y(n9361) );
  MUX2X1 U10916 ( .B(ram[2371]), .A(ram[2387]), .S(n12625), .Y(n9360) );
  MUX2X1 U10917 ( .B(ram[2339]), .A(ram[2355]), .S(n12632), .Y(n9364) );
  MUX2X1 U10918 ( .B(ram[2307]), .A(ram[2323]), .S(n12640), .Y(n9363) );
  MUX2X1 U10919 ( .B(n9362), .A(n9359), .S(mem_access_addr[2]), .Y(n9366) );
  MUX2X1 U10920 ( .B(ram[2275]), .A(ram[2291]), .S(n12662), .Y(n9370) );
  MUX2X1 U10921 ( .B(ram[2243]), .A(ram[2259]), .S(n12661), .Y(n9369) );
  MUX2X1 U10922 ( .B(ram[2211]), .A(ram[2227]), .S(n12621), .Y(n9373) );
  MUX2X1 U10923 ( .B(ram[2179]), .A(ram[2195]), .S(n12673), .Y(n9372) );
  MUX2X1 U10924 ( .B(n9371), .A(n9368), .S(n12587), .Y(n9382) );
  MUX2X1 U10925 ( .B(ram[2147]), .A(ram[2163]), .S(n12659), .Y(n9376) );
  MUX2X1 U10926 ( .B(ram[2115]), .A(ram[2131]), .S(n12621), .Y(n9375) );
  MUX2X1 U10927 ( .B(ram[2083]), .A(ram[2099]), .S(n12631), .Y(n9379) );
  MUX2X1 U10928 ( .B(ram[2051]), .A(ram[2067]), .S(n12642), .Y(n9378) );
  MUX2X1 U10929 ( .B(n9377), .A(n9374), .S(n12587), .Y(n9381) );
  MUX2X1 U10930 ( .B(n9380), .A(n9365), .S(n12564), .Y(n9384) );
  MUX2X1 U10931 ( .B(n9383), .A(n9320), .S(mem_access_addr[6]), .Y(n9513) );
  MUX2X1 U10932 ( .B(ram[2019]), .A(ram[2035]), .S(n12633), .Y(n9388) );
  MUX2X1 U10933 ( .B(ram[1987]), .A(ram[2003]), .S(n12675), .Y(n9387) );
  MUX2X1 U10934 ( .B(ram[1955]), .A(ram[1971]), .S(n12651), .Y(n9391) );
  MUX2X1 U10935 ( .B(ram[1923]), .A(ram[1939]), .S(n12673), .Y(n9390) );
  MUX2X1 U10936 ( .B(n9389), .A(n9386), .S(n12582), .Y(n9400) );
  MUX2X1 U10937 ( .B(ram[1891]), .A(ram[1907]), .S(n12648), .Y(n9394) );
  MUX2X1 U10938 ( .B(ram[1859]), .A(ram[1875]), .S(n12637), .Y(n9393) );
  MUX2X1 U10939 ( .B(ram[1827]), .A(ram[1843]), .S(n12682), .Y(n9397) );
  MUX2X1 U10940 ( .B(ram[1795]), .A(ram[1811]), .S(n12668), .Y(n9396) );
  MUX2X1 U10941 ( .B(n9395), .A(n9392), .S(n12582), .Y(n9399) );
  MUX2X1 U10942 ( .B(ram[1763]), .A(ram[1779]), .S(n12671), .Y(n9403) );
  MUX2X1 U10943 ( .B(ram[1731]), .A(ram[1747]), .S(n12669), .Y(n9402) );
  MUX2X1 U10944 ( .B(ram[1699]), .A(ram[1715]), .S(n12676), .Y(n9406) );
  MUX2X1 U10945 ( .B(ram[1667]), .A(ram[1683]), .S(n12634), .Y(n9405) );
  MUX2X1 U10946 ( .B(n9404), .A(n9401), .S(n12584), .Y(n9415) );
  MUX2X1 U10947 ( .B(ram[1635]), .A(ram[1651]), .S(n12659), .Y(n9409) );
  MUX2X1 U10948 ( .B(ram[1603]), .A(ram[1619]), .S(n12628), .Y(n9408) );
  MUX2X1 U10949 ( .B(ram[1571]), .A(ram[1587]), .S(n12679), .Y(n9412) );
  MUX2X1 U10950 ( .B(ram[1539]), .A(ram[1555]), .S(n12679), .Y(n9411) );
  MUX2X1 U10951 ( .B(n9410), .A(n9407), .S(mem_access_addr[2]), .Y(n9414) );
  MUX2X1 U10952 ( .B(n9413), .A(n9398), .S(n12566), .Y(n9448) );
  MUX2X1 U10953 ( .B(ram[1507]), .A(ram[1523]), .S(n12649), .Y(n9418) );
  MUX2X1 U10954 ( .B(ram[1475]), .A(ram[1491]), .S(n12681), .Y(n9417) );
  MUX2X1 U10955 ( .B(ram[1443]), .A(ram[1459]), .S(n12654), .Y(n9421) );
  MUX2X1 U10956 ( .B(ram[1411]), .A(ram[1427]), .S(n12647), .Y(n9420) );
  MUX2X1 U10957 ( .B(n9419), .A(n9416), .S(n12588), .Y(n9430) );
  MUX2X1 U10958 ( .B(ram[1379]), .A(ram[1395]), .S(n12631), .Y(n9424) );
  MUX2X1 U10959 ( .B(ram[1347]), .A(ram[1363]), .S(n12655), .Y(n9423) );
  MUX2X1 U10960 ( .B(ram[1315]), .A(ram[1331]), .S(n12643), .Y(n9427) );
  MUX2X1 U10961 ( .B(ram[1283]), .A(ram[1299]), .S(n12637), .Y(n9426) );
  MUX2X1 U10962 ( .B(n9425), .A(n9422), .S(n12581), .Y(n9429) );
  MUX2X1 U10963 ( .B(ram[1251]), .A(ram[1267]), .S(n12630), .Y(n9433) );
  MUX2X1 U10964 ( .B(ram[1219]), .A(ram[1235]), .S(n12670), .Y(n9432) );
  MUX2X1 U10965 ( .B(ram[1187]), .A(ram[1203]), .S(n12676), .Y(n9436) );
  MUX2X1 U10966 ( .B(ram[1155]), .A(ram[1171]), .S(n12657), .Y(n9435) );
  MUX2X1 U10967 ( .B(n9434), .A(n9431), .S(n12584), .Y(n9445) );
  MUX2X1 U10968 ( .B(ram[1123]), .A(ram[1139]), .S(n12649), .Y(n9439) );
  MUX2X1 U10969 ( .B(ram[1091]), .A(ram[1107]), .S(n12678), .Y(n9438) );
  MUX2X1 U10970 ( .B(ram[1059]), .A(ram[1075]), .S(n12666), .Y(n9442) );
  MUX2X1 U10971 ( .B(ram[1027]), .A(ram[1043]), .S(n12681), .Y(n9441) );
  MUX2X1 U10972 ( .B(n9440), .A(n9437), .S(n12582), .Y(n9444) );
  MUX2X1 U10973 ( .B(n9443), .A(n9428), .S(n12564), .Y(n9447) );
  MUX2X1 U10974 ( .B(ram[995]), .A(ram[1011]), .S(n12672), .Y(n9451) );
  MUX2X1 U10975 ( .B(ram[963]), .A(ram[979]), .S(n12640), .Y(n9450) );
  MUX2X1 U10976 ( .B(ram[931]), .A(ram[947]), .S(n12677), .Y(n9454) );
  MUX2X1 U10977 ( .B(ram[899]), .A(ram[915]), .S(n12657), .Y(n9453) );
  MUX2X1 U10978 ( .B(n9452), .A(n9449), .S(n12588), .Y(n9463) );
  MUX2X1 U10979 ( .B(ram[867]), .A(ram[883]), .S(n12676), .Y(n9457) );
  MUX2X1 U10980 ( .B(ram[835]), .A(ram[851]), .S(n12669), .Y(n9456) );
  MUX2X1 U10981 ( .B(ram[803]), .A(ram[819]), .S(n12655), .Y(n9460) );
  MUX2X1 U10982 ( .B(ram[771]), .A(ram[787]), .S(n12623), .Y(n9459) );
  MUX2X1 U10983 ( .B(n9458), .A(n9455), .S(n12576), .Y(n9462) );
  MUX2X1 U10984 ( .B(ram[739]), .A(ram[755]), .S(n12638), .Y(n9466) );
  MUX2X1 U10985 ( .B(ram[707]), .A(ram[723]), .S(n12667), .Y(n9465) );
  MUX2X1 U10986 ( .B(ram[675]), .A(ram[691]), .S(n12621), .Y(n9469) );
  MUX2X1 U10987 ( .B(ram[643]), .A(ram[659]), .S(n12676), .Y(n9468) );
  MUX2X1 U10988 ( .B(n9467), .A(n9464), .S(n12583), .Y(n9478) );
  MUX2X1 U10989 ( .B(ram[611]), .A(ram[627]), .S(n12630), .Y(n9472) );
  MUX2X1 U10990 ( .B(ram[579]), .A(ram[595]), .S(n12657), .Y(n9471) );
  MUX2X1 U10991 ( .B(ram[547]), .A(ram[563]), .S(n12656), .Y(n9475) );
  MUX2X1 U10992 ( .B(ram[515]), .A(ram[531]), .S(mem_access_addr[0]), .Y(n9474) );
  MUX2X1 U10993 ( .B(n9473), .A(n9470), .S(n12580), .Y(n9477) );
  MUX2X1 U10994 ( .B(n9476), .A(n9461), .S(n12566), .Y(n9511) );
  MUX2X1 U10995 ( .B(ram[483]), .A(ram[499]), .S(n12644), .Y(n9481) );
  MUX2X1 U10996 ( .B(ram[451]), .A(ram[467]), .S(n12660), .Y(n9480) );
  MUX2X1 U10997 ( .B(ram[419]), .A(ram[435]), .S(n12673), .Y(n9484) );
  MUX2X1 U10998 ( .B(ram[387]), .A(ram[403]), .S(mem_access_addr[0]), .Y(n9483) );
  MUX2X1 U10999 ( .B(n9482), .A(n9479), .S(n12576), .Y(n9493) );
  MUX2X1 U11000 ( .B(ram[355]), .A(ram[371]), .S(n12659), .Y(n9487) );
  MUX2X1 U11001 ( .B(ram[323]), .A(ram[339]), .S(n12634), .Y(n9486) );
  MUX2X1 U11002 ( .B(ram[291]), .A(ram[307]), .S(n12621), .Y(n9490) );
  MUX2X1 U11003 ( .B(ram[259]), .A(ram[275]), .S(mem_access_addr[0]), .Y(n9489) );
  MUX2X1 U11004 ( .B(n9488), .A(n9485), .S(n12580), .Y(n9492) );
  MUX2X1 U11005 ( .B(ram[227]), .A(ram[243]), .S(n12672), .Y(n9496) );
  MUX2X1 U11006 ( .B(ram[195]), .A(ram[211]), .S(n12671), .Y(n9495) );
  MUX2X1 U11007 ( .B(ram[163]), .A(ram[179]), .S(n12681), .Y(n9499) );
  MUX2X1 U11008 ( .B(ram[131]), .A(ram[147]), .S(n12633), .Y(n9498) );
  MUX2X1 U11009 ( .B(n9497), .A(n9494), .S(n12575), .Y(n9508) );
  MUX2X1 U11010 ( .B(ram[99]), .A(ram[115]), .S(n12661), .Y(n9502) );
  MUX2X1 U11011 ( .B(ram[67]), .A(ram[83]), .S(n12648), .Y(n9501) );
  MUX2X1 U11012 ( .B(ram[35]), .A(ram[51]), .S(mem_access_addr[0]), .Y(n9505)
         );
  MUX2X1 U11013 ( .B(ram[3]), .A(ram[19]), .S(n12658), .Y(n9504) );
  MUX2X1 U11014 ( .B(n9503), .A(n9500), .S(n12579), .Y(n9507) );
  MUX2X1 U11015 ( .B(n9506), .A(n9491), .S(n12567), .Y(n9510) );
  MUX2X1 U11016 ( .B(n9509), .A(n9446), .S(mem_access_addr[6]), .Y(n9512) );
  MUX2X1 U11017 ( .B(ram[4068]), .A(ram[4084]), .S(n12625), .Y(n9516) );
  MUX2X1 U11018 ( .B(ram[4036]), .A(ram[4052]), .S(n12628), .Y(n9515) );
  MUX2X1 U11019 ( .B(ram[4004]), .A(ram[4020]), .S(n12632), .Y(n9519) );
  MUX2X1 U11020 ( .B(ram[3972]), .A(ram[3988]), .S(n12626), .Y(n9518) );
  MUX2X1 U11021 ( .B(n9517), .A(n9514), .S(n12584), .Y(n9528) );
  MUX2X1 U11022 ( .B(ram[3940]), .A(ram[3956]), .S(n12630), .Y(n9522) );
  MUX2X1 U11023 ( .B(ram[3908]), .A(ram[3924]), .S(n12641), .Y(n9521) );
  MUX2X1 U11024 ( .B(ram[3876]), .A(ram[3892]), .S(n12633), .Y(n9525) );
  MUX2X1 U11025 ( .B(ram[3844]), .A(ram[3860]), .S(n12682), .Y(n9524) );
  MUX2X1 U11026 ( .B(n9523), .A(n9520), .S(n12583), .Y(n9527) );
  MUX2X1 U11027 ( .B(ram[3812]), .A(ram[3828]), .S(n12657), .Y(n9531) );
  MUX2X1 U11028 ( .B(ram[3780]), .A(ram[3796]), .S(n12629), .Y(n9530) );
  MUX2X1 U11029 ( .B(ram[3748]), .A(ram[3764]), .S(n12680), .Y(n9534) );
  MUX2X1 U11030 ( .B(ram[3716]), .A(ram[3732]), .S(n12667), .Y(n9533) );
  MUX2X1 U11031 ( .B(n9532), .A(n9529), .S(n12588), .Y(n9543) );
  MUX2X1 U11032 ( .B(ram[3684]), .A(ram[3700]), .S(n12623), .Y(n9537) );
  MUX2X1 U11033 ( .B(ram[3652]), .A(ram[3668]), .S(n12634), .Y(n9536) );
  MUX2X1 U11034 ( .B(ram[3620]), .A(ram[3636]), .S(n12635), .Y(n9540) );
  MUX2X1 U11035 ( .B(ram[3588]), .A(ram[3604]), .S(n12633), .Y(n9539) );
  MUX2X1 U11036 ( .B(n9538), .A(n9535), .S(n12577), .Y(n9542) );
  MUX2X1 U11037 ( .B(n9541), .A(n9526), .S(n12567), .Y(n9576) );
  MUX2X1 U11038 ( .B(ram[3556]), .A(ram[3572]), .S(mem_access_addr[0]), .Y(
        n9546) );
  MUX2X1 U11039 ( .B(ram[3524]), .A(ram[3540]), .S(n12622), .Y(n9545) );
  MUX2X1 U11040 ( .B(ram[3492]), .A(ram[3508]), .S(n12625), .Y(n9549) );
  MUX2X1 U11041 ( .B(ram[3460]), .A(ram[3476]), .S(n12653), .Y(n9548) );
  MUX2X1 U11042 ( .B(n9547), .A(n9544), .S(n12581), .Y(n9558) );
  MUX2X1 U11043 ( .B(ram[3428]), .A(ram[3444]), .S(n12637), .Y(n9552) );
  MUX2X1 U11044 ( .B(ram[3396]), .A(ram[3412]), .S(n12651), .Y(n9551) );
  MUX2X1 U11045 ( .B(ram[3364]), .A(ram[3380]), .S(n12666), .Y(n9555) );
  MUX2X1 U11046 ( .B(ram[3332]), .A(ram[3348]), .S(n12662), .Y(n9554) );
  MUX2X1 U11047 ( .B(n9553), .A(n9550), .S(n12589), .Y(n9557) );
  MUX2X1 U11048 ( .B(ram[3300]), .A(ram[3316]), .S(n12628), .Y(n9561) );
  MUX2X1 U11049 ( .B(ram[3268]), .A(ram[3284]), .S(n12636), .Y(n9560) );
  MUX2X1 U11050 ( .B(ram[3236]), .A(ram[3252]), .S(n12626), .Y(n9564) );
  MUX2X1 U11051 ( .B(ram[3204]), .A(ram[3220]), .S(n12673), .Y(n9563) );
  MUX2X1 U11052 ( .B(n9562), .A(n9559), .S(n12586), .Y(n9573) );
  MUX2X1 U11053 ( .B(ram[3172]), .A(ram[3188]), .S(n12628), .Y(n9567) );
  MUX2X1 U11054 ( .B(ram[3140]), .A(ram[3156]), .S(n12675), .Y(n9566) );
  MUX2X1 U11055 ( .B(ram[3108]), .A(ram[3124]), .S(n12636), .Y(n9570) );
  MUX2X1 U11056 ( .B(ram[3076]), .A(ram[3092]), .S(n12658), .Y(n9569) );
  MUX2X1 U11057 ( .B(n9568), .A(n9565), .S(n12582), .Y(n9572) );
  MUX2X1 U11058 ( .B(n9571), .A(n9556), .S(n12567), .Y(n9575) );
  MUX2X1 U11059 ( .B(ram[3044]), .A(ram[3060]), .S(n12627), .Y(n9579) );
  MUX2X1 U11060 ( .B(ram[3012]), .A(ram[3028]), .S(n12633), .Y(n9578) );
  MUX2X1 U11061 ( .B(ram[2980]), .A(ram[2996]), .S(n12648), .Y(n9582) );
  MUX2X1 U11062 ( .B(ram[2948]), .A(ram[2964]), .S(n12650), .Y(n9581) );
  MUX2X1 U11063 ( .B(n9580), .A(n9577), .S(n12575), .Y(n9591) );
  MUX2X1 U11064 ( .B(ram[2916]), .A(ram[2932]), .S(n12634), .Y(n9585) );
  MUX2X1 U11065 ( .B(ram[2884]), .A(ram[2900]), .S(n12629), .Y(n9584) );
  MUX2X1 U11066 ( .B(ram[2852]), .A(ram[2868]), .S(n12622), .Y(n9588) );
  MUX2X1 U11067 ( .B(ram[2820]), .A(ram[2836]), .S(n12643), .Y(n9587) );
  MUX2X1 U11068 ( .B(n9586), .A(n9583), .S(n12580), .Y(n9590) );
  MUX2X1 U11069 ( .B(ram[2788]), .A(ram[2804]), .S(n12631), .Y(n9594) );
  MUX2X1 U11070 ( .B(ram[2756]), .A(ram[2772]), .S(n12638), .Y(n9593) );
  MUX2X1 U11071 ( .B(ram[2724]), .A(ram[2740]), .S(n12636), .Y(n9597) );
  MUX2X1 U11072 ( .B(ram[2692]), .A(ram[2708]), .S(n12630), .Y(n9596) );
  MUX2X1 U11073 ( .B(n9595), .A(n9592), .S(n12575), .Y(n9606) );
  MUX2X1 U11074 ( .B(ram[2660]), .A(ram[2676]), .S(n12657), .Y(n9600) );
  MUX2X1 U11075 ( .B(ram[2628]), .A(ram[2644]), .S(n12644), .Y(n9599) );
  MUX2X1 U11076 ( .B(ram[2596]), .A(ram[2612]), .S(n12625), .Y(n9603) );
  MUX2X1 U11077 ( .B(ram[2564]), .A(ram[2580]), .S(n12633), .Y(n9602) );
  MUX2X1 U11078 ( .B(n9601), .A(n9598), .S(n12588), .Y(n9605) );
  MUX2X1 U11079 ( .B(n9604), .A(n9589), .S(n12566), .Y(n9639) );
  MUX2X1 U11080 ( .B(ram[2532]), .A(ram[2548]), .S(n12674), .Y(n9609) );
  MUX2X1 U11081 ( .B(ram[2500]), .A(ram[2516]), .S(n12648), .Y(n9608) );
  MUX2X1 U11082 ( .B(ram[2468]), .A(ram[2484]), .S(n12634), .Y(n9612) );
  MUX2X1 U11083 ( .B(ram[2436]), .A(ram[2452]), .S(n12661), .Y(n9611) );
  MUX2X1 U11084 ( .B(n9610), .A(n9607), .S(n12584), .Y(n9621) );
  MUX2X1 U11085 ( .B(ram[2404]), .A(ram[2420]), .S(n12661), .Y(n9615) );
  MUX2X1 U11086 ( .B(ram[2372]), .A(ram[2388]), .S(n12658), .Y(n9614) );
  MUX2X1 U11087 ( .B(ram[2340]), .A(ram[2356]), .S(n12674), .Y(n9618) );
  MUX2X1 U11088 ( .B(ram[2308]), .A(ram[2324]), .S(n12627), .Y(n9617) );
  MUX2X1 U11089 ( .B(n9616), .A(n9613), .S(n12588), .Y(n9620) );
  MUX2X1 U11090 ( .B(ram[2276]), .A(ram[2292]), .S(n12626), .Y(n9624) );
  MUX2X1 U11091 ( .B(ram[2244]), .A(ram[2260]), .S(n12635), .Y(n9623) );
  MUX2X1 U11092 ( .B(ram[2212]), .A(ram[2228]), .S(n12637), .Y(n9627) );
  MUX2X1 U11093 ( .B(ram[2180]), .A(ram[2196]), .S(n12642), .Y(n9626) );
  MUX2X1 U11094 ( .B(n9625), .A(n9622), .S(n12579), .Y(n9636) );
  MUX2X1 U11095 ( .B(ram[2148]), .A(ram[2164]), .S(n12680), .Y(n9630) );
  MUX2X1 U11096 ( .B(ram[2116]), .A(ram[2132]), .S(n12660), .Y(n9629) );
  MUX2X1 U11097 ( .B(ram[2084]), .A(ram[2100]), .S(n12627), .Y(n9633) );
  MUX2X1 U11098 ( .B(ram[2052]), .A(ram[2068]), .S(n12638), .Y(n9632) );
  MUX2X1 U11099 ( .B(n9631), .A(n9628), .S(n12588), .Y(n9635) );
  MUX2X1 U11100 ( .B(n9634), .A(n9619), .S(n12565), .Y(n9638) );
  MUX2X1 U11101 ( .B(n9637), .A(n9574), .S(mem_access_addr[6]), .Y(n9767) );
  MUX2X1 U11102 ( .B(ram[2020]), .A(ram[2036]), .S(n12648), .Y(n9642) );
  MUX2X1 U11103 ( .B(ram[1988]), .A(ram[2004]), .S(n12665), .Y(n9641) );
  MUX2X1 U11104 ( .B(ram[1956]), .A(ram[1972]), .S(n12630), .Y(n9645) );
  MUX2X1 U11105 ( .B(ram[1924]), .A(ram[1940]), .S(n12665), .Y(n9644) );
  MUX2X1 U11106 ( .B(n9643), .A(n9640), .S(n12589), .Y(n9654) );
  MUX2X1 U11107 ( .B(ram[1892]), .A(ram[1908]), .S(n12675), .Y(n9648) );
  MUX2X1 U11108 ( .B(ram[1860]), .A(ram[1876]), .S(n12646), .Y(n9647) );
  MUX2X1 U11109 ( .B(ram[1828]), .A(ram[1844]), .S(n12630), .Y(n9651) );
  MUX2X1 U11110 ( .B(ram[1796]), .A(ram[1812]), .S(n12676), .Y(n9650) );
  MUX2X1 U11111 ( .B(n9649), .A(n9646), .S(n12586), .Y(n9653) );
  MUX2X1 U11112 ( .B(ram[1764]), .A(ram[1780]), .S(n12674), .Y(n9657) );
  MUX2X1 U11113 ( .B(ram[1732]), .A(ram[1748]), .S(n12655), .Y(n9656) );
  MUX2X1 U11114 ( .B(ram[1700]), .A(ram[1716]), .S(n12634), .Y(n9660) );
  MUX2X1 U11115 ( .B(ram[1668]), .A(ram[1684]), .S(n12683), .Y(n9659) );
  MUX2X1 U11116 ( .B(n9658), .A(n9655), .S(n12589), .Y(n9669) );
  MUX2X1 U11117 ( .B(ram[1636]), .A(ram[1652]), .S(n12624), .Y(n9663) );
  MUX2X1 U11118 ( .B(ram[1604]), .A(ram[1620]), .S(n12638), .Y(n9662) );
  MUX2X1 U11119 ( .B(ram[1572]), .A(ram[1588]), .S(n12656), .Y(n9666) );
  MUX2X1 U11120 ( .B(ram[1540]), .A(ram[1556]), .S(n12622), .Y(n9665) );
  MUX2X1 U11121 ( .B(n9664), .A(n9661), .S(n12587), .Y(n9668) );
  MUX2X1 U11122 ( .B(n9667), .A(n9652), .S(n12566), .Y(n9702) );
  MUX2X1 U11123 ( .B(ram[1508]), .A(ram[1524]), .S(n12649), .Y(n9672) );
  MUX2X1 U11124 ( .B(ram[1476]), .A(ram[1492]), .S(n12651), .Y(n9671) );
  MUX2X1 U11125 ( .B(ram[1444]), .A(ram[1460]), .S(n12623), .Y(n9675) );
  MUX2X1 U11126 ( .B(ram[1412]), .A(ram[1428]), .S(n12641), .Y(n9674) );
  MUX2X1 U11127 ( .B(n9673), .A(n9670), .S(n12587), .Y(n9684) );
  MUX2X1 U11128 ( .B(ram[1380]), .A(ram[1396]), .S(n12634), .Y(n9678) );
  MUX2X1 U11129 ( .B(ram[1348]), .A(ram[1364]), .S(n12664), .Y(n9677) );
  MUX2X1 U11130 ( .B(ram[1316]), .A(ram[1332]), .S(n12682), .Y(n9681) );
  MUX2X1 U11131 ( .B(ram[1284]), .A(ram[1300]), .S(n12661), .Y(n9680) );
  MUX2X1 U11132 ( .B(n9679), .A(n9676), .S(n12587), .Y(n9683) );
  MUX2X1 U11133 ( .B(ram[1252]), .A(ram[1268]), .S(mem_access_addr[0]), .Y(
        n9687) );
  MUX2X1 U11134 ( .B(ram[1220]), .A(ram[1236]), .S(n12668), .Y(n9686) );
  MUX2X1 U11135 ( .B(ram[1188]), .A(ram[1204]), .S(n12659), .Y(n9690) );
  MUX2X1 U11136 ( .B(ram[1156]), .A(ram[1172]), .S(n12677), .Y(n9689) );
  MUX2X1 U11137 ( .B(n9688), .A(n9685), .S(n12586), .Y(n9699) );
  MUX2X1 U11138 ( .B(ram[1124]), .A(ram[1140]), .S(n12649), .Y(n9693) );
  MUX2X1 U11139 ( .B(ram[1092]), .A(ram[1108]), .S(n12663), .Y(n9692) );
  MUX2X1 U11140 ( .B(ram[1060]), .A(ram[1076]), .S(n12675), .Y(n9696) );
  MUX2X1 U11141 ( .B(ram[1028]), .A(ram[1044]), .S(n12638), .Y(n9695) );
  MUX2X1 U11142 ( .B(n9694), .A(n9691), .S(n12580), .Y(n9698) );
  MUX2X1 U11143 ( .B(n9697), .A(n9682), .S(n12565), .Y(n9701) );
  MUX2X1 U11144 ( .B(ram[996]), .A(ram[1012]), .S(n12638), .Y(n9705) );
  MUX2X1 U11145 ( .B(ram[964]), .A(ram[980]), .S(n12681), .Y(n9704) );
  MUX2X1 U11146 ( .B(ram[932]), .A(ram[948]), .S(n12631), .Y(n9708) );
  MUX2X1 U11147 ( .B(ram[900]), .A(ram[916]), .S(n12627), .Y(n9707) );
  MUX2X1 U11148 ( .B(n9706), .A(n9703), .S(n12587), .Y(n9717) );
  MUX2X1 U11149 ( .B(ram[868]), .A(ram[884]), .S(n12656), .Y(n9711) );
  MUX2X1 U11150 ( .B(ram[836]), .A(ram[852]), .S(n12621), .Y(n9710) );
  MUX2X1 U11151 ( .B(ram[804]), .A(ram[820]), .S(n12639), .Y(n9714) );
  MUX2X1 U11152 ( .B(ram[772]), .A(ram[788]), .S(n12659), .Y(n9713) );
  MUX2X1 U11153 ( .B(n9712), .A(n9709), .S(n12585), .Y(n9716) );
  MUX2X1 U11154 ( .B(ram[740]), .A(ram[756]), .S(n12632), .Y(n9720) );
  MUX2X1 U11155 ( .B(ram[708]), .A(ram[724]), .S(n12640), .Y(n9719) );
  MUX2X1 U11156 ( .B(ram[676]), .A(ram[692]), .S(n12625), .Y(n9723) );
  MUX2X1 U11157 ( .B(ram[644]), .A(ram[660]), .S(n12670), .Y(n9722) );
  MUX2X1 U11158 ( .B(n9721), .A(n9718), .S(n12589), .Y(n9732) );
  MUX2X1 U11159 ( .B(ram[612]), .A(ram[628]), .S(n12636), .Y(n9726) );
  MUX2X1 U11160 ( .B(ram[580]), .A(ram[596]), .S(n12678), .Y(n9725) );
  MUX2X1 U11161 ( .B(ram[548]), .A(ram[564]), .S(n12656), .Y(n9729) );
  MUX2X1 U11162 ( .B(ram[516]), .A(ram[532]), .S(n12632), .Y(n9728) );
  MUX2X1 U11163 ( .B(n9727), .A(n9724), .S(n12586), .Y(n9731) );
  MUX2X1 U11164 ( .B(n9730), .A(n9715), .S(n12567), .Y(n9765) );
  MUX2X1 U11165 ( .B(ram[484]), .A(ram[500]), .S(n12641), .Y(n9735) );
  MUX2X1 U11166 ( .B(ram[452]), .A(ram[468]), .S(n12645), .Y(n9734) );
  MUX2X1 U11167 ( .B(ram[420]), .A(ram[436]), .S(n12662), .Y(n9738) );
  MUX2X1 U11168 ( .B(ram[388]), .A(ram[404]), .S(n12643), .Y(n9737) );
  MUX2X1 U11169 ( .B(n9736), .A(n9733), .S(n12586), .Y(n9747) );
  MUX2X1 U11170 ( .B(ram[356]), .A(ram[372]), .S(n12647), .Y(n9741) );
  MUX2X1 U11171 ( .B(ram[324]), .A(ram[340]), .S(n12657), .Y(n9740) );
  MUX2X1 U11172 ( .B(ram[292]), .A(ram[308]), .S(n12644), .Y(n9744) );
  MUX2X1 U11173 ( .B(ram[260]), .A(ram[276]), .S(n12631), .Y(n9743) );
  MUX2X1 U11174 ( .B(n9742), .A(n9739), .S(n12586), .Y(n9746) );
  MUX2X1 U11175 ( .B(ram[228]), .A(ram[244]), .S(n12638), .Y(n9750) );
  MUX2X1 U11176 ( .B(ram[196]), .A(ram[212]), .S(n12643), .Y(n9749) );
  MUX2X1 U11177 ( .B(ram[164]), .A(ram[180]), .S(n12678), .Y(n9753) );
  MUX2X1 U11178 ( .B(ram[132]), .A(ram[148]), .S(n12627), .Y(n9752) );
  MUX2X1 U11179 ( .B(n9751), .A(n9748), .S(n12589), .Y(n9762) );
  MUX2X1 U11180 ( .B(ram[100]), .A(ram[116]), .S(mem_access_addr[0]), .Y(n9756) );
  MUX2X1 U11181 ( .B(ram[68]), .A(ram[84]), .S(n12643), .Y(n9755) );
  MUX2X1 U11182 ( .B(ram[36]), .A(ram[52]), .S(n12626), .Y(n9759) );
  MUX2X1 U11183 ( .B(ram[4]), .A(ram[20]), .S(n12646), .Y(n9758) );
  MUX2X1 U11184 ( .B(n9757), .A(n9754), .S(n12586), .Y(n9761) );
  MUX2X1 U11185 ( .B(n9760), .A(n9745), .S(n12566), .Y(n9764) );
  MUX2X1 U11186 ( .B(n9763), .A(n9700), .S(mem_access_addr[6]), .Y(n9766) );
  MUX2X1 U11187 ( .B(ram[4069]), .A(ram[4085]), .S(n12623), .Y(n9770) );
  MUX2X1 U11188 ( .B(ram[4037]), .A(ram[4053]), .S(n12663), .Y(n9769) );
  MUX2X1 U11189 ( .B(ram[4005]), .A(ram[4021]), .S(n12647), .Y(n9773) );
  MUX2X1 U11190 ( .B(ram[3973]), .A(ram[3989]), .S(n12649), .Y(n9772) );
  MUX2X1 U11191 ( .B(n9771), .A(n9768), .S(n12579), .Y(n9782) );
  MUX2X1 U11192 ( .B(ram[3941]), .A(ram[3957]), .S(n12660), .Y(n9776) );
  MUX2X1 U11193 ( .B(ram[3909]), .A(ram[3925]), .S(n12633), .Y(n9775) );
  MUX2X1 U11194 ( .B(ram[3877]), .A(ram[3893]), .S(n12660), .Y(n9779) );
  MUX2X1 U11195 ( .B(ram[3845]), .A(ram[3861]), .S(n12657), .Y(n9778) );
  MUX2X1 U11196 ( .B(n9777), .A(n9774), .S(n12586), .Y(n9781) );
  MUX2X1 U11197 ( .B(ram[3813]), .A(ram[3829]), .S(n12674), .Y(n9785) );
  MUX2X1 U11198 ( .B(ram[3781]), .A(ram[3797]), .S(n12675), .Y(n9784) );
  MUX2X1 U11199 ( .B(ram[3749]), .A(ram[3765]), .S(n12627), .Y(n9788) );
  MUX2X1 U11200 ( .B(ram[3717]), .A(ram[3733]), .S(n12628), .Y(n9787) );
  MUX2X1 U11201 ( .B(n9786), .A(n9783), .S(n12588), .Y(n9797) );
  MUX2X1 U11202 ( .B(ram[3685]), .A(ram[3701]), .S(n12646), .Y(n9791) );
  MUX2X1 U11203 ( .B(ram[3653]), .A(ram[3669]), .S(n12658), .Y(n9790) );
  MUX2X1 U11204 ( .B(ram[3621]), .A(ram[3637]), .S(n12635), .Y(n9794) );
  MUX2X1 U11205 ( .B(ram[3589]), .A(ram[3605]), .S(n12667), .Y(n9793) );
  MUX2X1 U11206 ( .B(n9792), .A(n9789), .S(n12585), .Y(n9796) );
  MUX2X1 U11207 ( .B(n9795), .A(n9780), .S(n12564), .Y(n9830) );
  MUX2X1 U11208 ( .B(ram[3557]), .A(ram[3573]), .S(n12638), .Y(n9800) );
  MUX2X1 U11209 ( .B(ram[3525]), .A(ram[3541]), .S(n12667), .Y(n9799) );
  MUX2X1 U11210 ( .B(ram[3493]), .A(ram[3509]), .S(n12649), .Y(n9803) );
  MUX2X1 U11211 ( .B(ram[3461]), .A(ram[3477]), .S(n12663), .Y(n9802) );
  MUX2X1 U11212 ( .B(n9801), .A(n9798), .S(n12586), .Y(n9812) );
  MUX2X1 U11213 ( .B(ram[3429]), .A(ram[3445]), .S(n12668), .Y(n9806) );
  MUX2X1 U11214 ( .B(ram[3397]), .A(ram[3413]), .S(n12641), .Y(n9805) );
  MUX2X1 U11215 ( .B(ram[3365]), .A(ram[3381]), .S(n12661), .Y(n9809) );
  MUX2X1 U11216 ( .B(ram[3333]), .A(ram[3349]), .S(n12627), .Y(n9808) );
  MUX2X1 U11217 ( .B(n9807), .A(n9804), .S(n12588), .Y(n9811) );
  MUX2X1 U11218 ( .B(ram[3301]), .A(ram[3317]), .S(n12682), .Y(n9815) );
  MUX2X1 U11219 ( .B(ram[3269]), .A(ram[3285]), .S(n12638), .Y(n9814) );
  MUX2X1 U11220 ( .B(ram[3237]), .A(ram[3253]), .S(n12630), .Y(n9818) );
  MUX2X1 U11221 ( .B(ram[3205]), .A(ram[3221]), .S(n12630), .Y(n9817) );
  MUX2X1 U11222 ( .B(n9816), .A(n9813), .S(n12585), .Y(n9827) );
  MUX2X1 U11223 ( .B(ram[3173]), .A(ram[3189]), .S(n12659), .Y(n9821) );
  MUX2X1 U11224 ( .B(ram[3141]), .A(ram[3157]), .S(n12627), .Y(n9820) );
  MUX2X1 U11225 ( .B(ram[3109]), .A(ram[3125]), .S(n12677), .Y(n9824) );
  MUX2X1 U11226 ( .B(ram[3077]), .A(ram[3093]), .S(n12656), .Y(n9823) );
  MUX2X1 U11227 ( .B(n9822), .A(n9819), .S(n12588), .Y(n9826) );
  MUX2X1 U11228 ( .B(n9825), .A(n9810), .S(n12565), .Y(n9829) );
  MUX2X1 U11229 ( .B(ram[3045]), .A(ram[3061]), .S(n12636), .Y(n9833) );
  MUX2X1 U11230 ( .B(ram[3013]), .A(ram[3029]), .S(n12662), .Y(n9832) );
  MUX2X1 U11231 ( .B(ram[2981]), .A(ram[2997]), .S(n12627), .Y(n9836) );
  MUX2X1 U11232 ( .B(ram[2949]), .A(ram[2965]), .S(n12676), .Y(n9835) );
  MUX2X1 U11233 ( .B(n9834), .A(n9831), .S(n12589), .Y(n9845) );
  MUX2X1 U11234 ( .B(ram[2917]), .A(ram[2933]), .S(n12673), .Y(n9839) );
  MUX2X1 U11235 ( .B(ram[2885]), .A(ram[2901]), .S(n12679), .Y(n9838) );
  MUX2X1 U11236 ( .B(ram[2853]), .A(ram[2869]), .S(n12642), .Y(n9842) );
  MUX2X1 U11237 ( .B(ram[2821]), .A(ram[2837]), .S(n12668), .Y(n9841) );
  MUX2X1 U11238 ( .B(n9840), .A(n9837), .S(n12580), .Y(n9844) );
  MUX2X1 U11239 ( .B(ram[2789]), .A(ram[2805]), .S(n12642), .Y(n9848) );
  MUX2X1 U11240 ( .B(ram[2757]), .A(ram[2773]), .S(n12664), .Y(n9847) );
  MUX2X1 U11241 ( .B(ram[2725]), .A(ram[2741]), .S(n12628), .Y(n9851) );
  MUX2X1 U11242 ( .B(ram[2693]), .A(ram[2709]), .S(n12631), .Y(n9850) );
  MUX2X1 U11243 ( .B(n9849), .A(n9846), .S(n12578), .Y(n9860) );
  MUX2X1 U11244 ( .B(ram[2661]), .A(ram[2677]), .S(n12666), .Y(n9854) );
  MUX2X1 U11245 ( .B(ram[2629]), .A(ram[2645]), .S(n12640), .Y(n9853) );
  MUX2X1 U11246 ( .B(ram[2597]), .A(ram[2613]), .S(n12637), .Y(n9857) );
  MUX2X1 U11247 ( .B(ram[2565]), .A(ram[2581]), .S(n12662), .Y(n9856) );
  MUX2X1 U11248 ( .B(n9855), .A(n9852), .S(n12584), .Y(n9859) );
  MUX2X1 U11249 ( .B(n9858), .A(n9843), .S(n12564), .Y(n9893) );
  MUX2X1 U11250 ( .B(ram[2533]), .A(ram[2549]), .S(n12670), .Y(n9863) );
  MUX2X1 U11251 ( .B(ram[2501]), .A(ram[2517]), .S(n12667), .Y(n9862) );
  MUX2X1 U11252 ( .B(ram[2469]), .A(ram[2485]), .S(n12653), .Y(n9866) );
  MUX2X1 U11253 ( .B(ram[2437]), .A(ram[2453]), .S(n12628), .Y(n9865) );
  MUX2X1 U11254 ( .B(n9864), .A(n9861), .S(n12576), .Y(n9875) );
  MUX2X1 U11255 ( .B(ram[2405]), .A(ram[2421]), .S(n12672), .Y(n9869) );
  MUX2X1 U11256 ( .B(ram[2373]), .A(ram[2389]), .S(n12657), .Y(n9868) );
  MUX2X1 U11257 ( .B(ram[2341]), .A(ram[2357]), .S(n12666), .Y(n9872) );
  MUX2X1 U11258 ( .B(ram[2309]), .A(ram[2325]), .S(n12652), .Y(n9871) );
  MUX2X1 U11259 ( .B(n9870), .A(n9867), .S(mem_access_addr[2]), .Y(n9874) );
  MUX2X1 U11260 ( .B(ram[2277]), .A(ram[2293]), .S(n12643), .Y(n9878) );
  MUX2X1 U11261 ( .B(ram[2245]), .A(ram[2261]), .S(n12665), .Y(n9877) );
  MUX2X1 U11262 ( .B(ram[2213]), .A(ram[2229]), .S(n12675), .Y(n9881) );
  MUX2X1 U11263 ( .B(ram[2181]), .A(ram[2197]), .S(n12630), .Y(n9880) );
  MUX2X1 U11264 ( .B(n9879), .A(n9876), .S(n12575), .Y(n9890) );
  MUX2X1 U11265 ( .B(ram[2149]), .A(ram[2165]), .S(n12650), .Y(n9884) );
  MUX2X1 U11266 ( .B(ram[2117]), .A(ram[2133]), .S(n12678), .Y(n9883) );
  MUX2X1 U11267 ( .B(ram[2085]), .A(ram[2101]), .S(n12654), .Y(n9887) );
  MUX2X1 U11268 ( .B(ram[2053]), .A(ram[2069]), .S(n12682), .Y(n9886) );
  MUX2X1 U11269 ( .B(n9885), .A(n9882), .S(n12578), .Y(n9889) );
  MUX2X1 U11270 ( .B(n9888), .A(n9873), .S(n12566), .Y(n9892) );
  MUX2X1 U11271 ( .B(n9891), .A(n9828), .S(mem_access_addr[6]), .Y(n10021) );
  MUX2X1 U11272 ( .B(ram[2021]), .A(ram[2037]), .S(n12643), .Y(n9896) );
  MUX2X1 U11273 ( .B(ram[1989]), .A(ram[2005]), .S(n12671), .Y(n9895) );
  MUX2X1 U11274 ( .B(ram[1957]), .A(ram[1973]), .S(n12654), .Y(n9899) );
  MUX2X1 U11275 ( .B(ram[1925]), .A(ram[1941]), .S(n12623), .Y(n9898) );
  MUX2X1 U11276 ( .B(n9897), .A(n9894), .S(n12586), .Y(n9908) );
  MUX2X1 U11277 ( .B(ram[1893]), .A(ram[1909]), .S(n12649), .Y(n9902) );
  MUX2X1 U11278 ( .B(ram[1861]), .A(ram[1877]), .S(n12663), .Y(n9901) );
  MUX2X1 U11279 ( .B(ram[1829]), .A(ram[1845]), .S(n12624), .Y(n9905) );
  MUX2X1 U11280 ( .B(ram[1797]), .A(ram[1813]), .S(n12654), .Y(n9904) );
  MUX2X1 U11281 ( .B(n9903), .A(n9900), .S(n12580), .Y(n9907) );
  MUX2X1 U11282 ( .B(ram[1765]), .A(ram[1781]), .S(n12648), .Y(n9911) );
  MUX2X1 U11283 ( .B(ram[1733]), .A(ram[1749]), .S(n12662), .Y(n9910) );
  MUX2X1 U11284 ( .B(ram[1701]), .A(ram[1717]), .S(n12644), .Y(n9914) );
  MUX2X1 U11285 ( .B(ram[1669]), .A(ram[1685]), .S(n12675), .Y(n9913) );
  MUX2X1 U11286 ( .B(n9912), .A(n9909), .S(n12580), .Y(n9923) );
  MUX2X1 U11287 ( .B(ram[1637]), .A(ram[1653]), .S(n12669), .Y(n9917) );
  MUX2X1 U11288 ( .B(ram[1605]), .A(ram[1621]), .S(n12624), .Y(n9916) );
  MUX2X1 U11289 ( .B(ram[1573]), .A(ram[1589]), .S(n12676), .Y(n9920) );
  MUX2X1 U11290 ( .B(ram[1541]), .A(ram[1557]), .S(n12663), .Y(n9919) );
  MUX2X1 U11291 ( .B(n9918), .A(n9915), .S(n12585), .Y(n9922) );
  MUX2X1 U11292 ( .B(n9921), .A(n9906), .S(n12566), .Y(n9956) );
  MUX2X1 U11293 ( .B(ram[1509]), .A(ram[1525]), .S(mem_access_addr[0]), .Y(
        n9926) );
  MUX2X1 U11294 ( .B(ram[1477]), .A(ram[1493]), .S(n12680), .Y(n9925) );
  MUX2X1 U11295 ( .B(ram[1445]), .A(ram[1461]), .S(n12661), .Y(n9929) );
  MUX2X1 U11296 ( .B(ram[1413]), .A(ram[1429]), .S(n12658), .Y(n9928) );
  MUX2X1 U11297 ( .B(n9927), .A(n9924), .S(n12583), .Y(n9938) );
  MUX2X1 U11298 ( .B(ram[1381]), .A(ram[1397]), .S(n12636), .Y(n9932) );
  MUX2X1 U11299 ( .B(ram[1349]), .A(ram[1365]), .S(n12657), .Y(n9931) );
  MUX2X1 U11300 ( .B(ram[1317]), .A(ram[1333]), .S(n12640), .Y(n9935) );
  MUX2X1 U11301 ( .B(ram[1285]), .A(ram[1301]), .S(n12648), .Y(n9934) );
  MUX2X1 U11302 ( .B(n9933), .A(n9930), .S(n12581), .Y(n9937) );
  MUX2X1 U11303 ( .B(ram[1253]), .A(ram[1269]), .S(n12679), .Y(n9941) );
  MUX2X1 U11304 ( .B(ram[1221]), .A(ram[1237]), .S(n12644), .Y(n9940) );
  MUX2X1 U11305 ( .B(ram[1189]), .A(ram[1205]), .S(n12673), .Y(n9944) );
  MUX2X1 U11306 ( .B(ram[1157]), .A(ram[1173]), .S(n12658), .Y(n9943) );
  MUX2X1 U11307 ( .B(n9942), .A(n9939), .S(n12579), .Y(n9953) );
  MUX2X1 U11308 ( .B(ram[1125]), .A(ram[1141]), .S(n12660), .Y(n9947) );
  MUX2X1 U11309 ( .B(ram[1093]), .A(ram[1109]), .S(n12675), .Y(n9946) );
  MUX2X1 U11310 ( .B(ram[1061]), .A(ram[1077]), .S(mem_access_addr[0]), .Y(
        n9950) );
  MUX2X1 U11311 ( .B(ram[1029]), .A(ram[1045]), .S(n12639), .Y(n9949) );
  MUX2X1 U11312 ( .B(n9948), .A(n9945), .S(n12577), .Y(n9952) );
  MUX2X1 U11313 ( .B(n9951), .A(n9936), .S(n12565), .Y(n9955) );
  MUX2X1 U11314 ( .B(ram[997]), .A(ram[1013]), .S(n12659), .Y(n9959) );
  MUX2X1 U11315 ( .B(ram[965]), .A(ram[981]), .S(n12656), .Y(n9958) );
  MUX2X1 U11316 ( .B(ram[933]), .A(ram[949]), .S(n12655), .Y(n9962) );
  MUX2X1 U11317 ( .B(ram[901]), .A(ram[917]), .S(n12677), .Y(n9961) );
  MUX2X1 U11318 ( .B(n9960), .A(n9957), .S(n12581), .Y(n9971) );
  MUX2X1 U11319 ( .B(ram[869]), .A(ram[885]), .S(n12645), .Y(n9965) );
  MUX2X1 U11320 ( .B(ram[837]), .A(ram[853]), .S(n12646), .Y(n9964) );
  MUX2X1 U11321 ( .B(ram[805]), .A(ram[821]), .S(n12632), .Y(n9968) );
  MUX2X1 U11322 ( .B(ram[773]), .A(ram[789]), .S(n12638), .Y(n9967) );
  MUX2X1 U11323 ( .B(n9966), .A(n9963), .S(n12587), .Y(n9970) );
  MUX2X1 U11324 ( .B(ram[741]), .A(ram[757]), .S(n12635), .Y(n9974) );
  MUX2X1 U11325 ( .B(ram[709]), .A(ram[725]), .S(n12622), .Y(n9973) );
  MUX2X1 U11326 ( .B(ram[677]), .A(ram[693]), .S(n12629), .Y(n9977) );
  MUX2X1 U11327 ( .B(ram[645]), .A(ram[661]), .S(n12637), .Y(n9976) );
  MUX2X1 U11328 ( .B(n9975), .A(n9972), .S(n12576), .Y(n9986) );
  MUX2X1 U11329 ( .B(ram[613]), .A(ram[629]), .S(n12624), .Y(n9980) );
  MUX2X1 U11330 ( .B(ram[581]), .A(ram[597]), .S(n12663), .Y(n9979) );
  MUX2X1 U11331 ( .B(ram[549]), .A(ram[565]), .S(n12632), .Y(n9983) );
  MUX2X1 U11332 ( .B(ram[517]), .A(ram[533]), .S(n12634), .Y(n9982) );
  MUX2X1 U11333 ( .B(n9981), .A(n9978), .S(n12580), .Y(n9985) );
  MUX2X1 U11334 ( .B(n9984), .A(n9969), .S(n12565), .Y(n10019) );
  MUX2X1 U11335 ( .B(ram[485]), .A(ram[501]), .S(n12662), .Y(n9989) );
  MUX2X1 U11336 ( .B(ram[453]), .A(ram[469]), .S(n12665), .Y(n9988) );
  MUX2X1 U11337 ( .B(ram[421]), .A(ram[437]), .S(n12679), .Y(n9992) );
  MUX2X1 U11338 ( .B(ram[389]), .A(ram[405]), .S(n12681), .Y(n9991) );
  MUX2X1 U11339 ( .B(n9990), .A(n9987), .S(mem_access_addr[2]), .Y(n10001) );
  MUX2X1 U11340 ( .B(ram[357]), .A(ram[373]), .S(n12637), .Y(n9995) );
  MUX2X1 U11341 ( .B(ram[325]), .A(ram[341]), .S(n12653), .Y(n9994) );
  MUX2X1 U11342 ( .B(ram[293]), .A(ram[309]), .S(n12646), .Y(n9998) );
  MUX2X1 U11343 ( .B(ram[261]), .A(ram[277]), .S(n12633), .Y(n9997) );
  MUX2X1 U11344 ( .B(n9996), .A(n9993), .S(mem_access_addr[2]), .Y(n10000) );
  MUX2X1 U11345 ( .B(ram[229]), .A(ram[245]), .S(n12623), .Y(n10004) );
  MUX2X1 U11346 ( .B(ram[197]), .A(ram[213]), .S(mem_access_addr[0]), .Y(
        n10003) );
  MUX2X1 U11347 ( .B(ram[165]), .A(ram[181]), .S(n12629), .Y(n10007) );
  MUX2X1 U11348 ( .B(ram[133]), .A(ram[149]), .S(n12624), .Y(n10006) );
  MUX2X1 U11349 ( .B(n10005), .A(n10002), .S(n12585), .Y(n10016) );
  MUX2X1 U11350 ( .B(ram[101]), .A(ram[117]), .S(n12654), .Y(n10010) );
  MUX2X1 U11351 ( .B(ram[69]), .A(ram[85]), .S(n12670), .Y(n10009) );
  MUX2X1 U11352 ( .B(ram[37]), .A(ram[53]), .S(n12633), .Y(n10013) );
  MUX2X1 U11353 ( .B(ram[5]), .A(ram[21]), .S(n12683), .Y(n10012) );
  MUX2X1 U11354 ( .B(n10011), .A(n10008), .S(mem_access_addr[2]), .Y(n10015)
         );
  MUX2X1 U11355 ( .B(n10014), .A(n9999), .S(n12565), .Y(n10018) );
  MUX2X1 U11356 ( .B(n10017), .A(n9954), .S(mem_access_addr[6]), .Y(n10020) );
  MUX2X1 U11357 ( .B(ram[4070]), .A(ram[4086]), .S(n12643), .Y(n10024) );
  MUX2X1 U11358 ( .B(ram[4038]), .A(ram[4054]), .S(n12669), .Y(n10023) );
  MUX2X1 U11359 ( .B(ram[4006]), .A(ram[4022]), .S(n12650), .Y(n10027) );
  MUX2X1 U11360 ( .B(ram[3974]), .A(ram[3990]), .S(n12682), .Y(n10026) );
  MUX2X1 U11361 ( .B(n10025), .A(n10022), .S(n12583), .Y(n10036) );
  MUX2X1 U11362 ( .B(ram[3942]), .A(ram[3958]), .S(n12641), .Y(n10030) );
  MUX2X1 U11363 ( .B(ram[3910]), .A(ram[3926]), .S(n12677), .Y(n10029) );
  MUX2X1 U11364 ( .B(ram[3878]), .A(ram[3894]), .S(n12652), .Y(n10033) );
  MUX2X1 U11365 ( .B(ram[3846]), .A(ram[3862]), .S(n12678), .Y(n10032) );
  MUX2X1 U11366 ( .B(n10031), .A(n10028), .S(mem_access_addr[2]), .Y(n10035)
         );
  MUX2X1 U11367 ( .B(ram[3814]), .A(ram[3830]), .S(n12632), .Y(n10039) );
  MUX2X1 U11368 ( .B(ram[3782]), .A(ram[3798]), .S(n12666), .Y(n10038) );
  MUX2X1 U11369 ( .B(ram[3750]), .A(ram[3766]), .S(n12644), .Y(n10042) );
  MUX2X1 U11370 ( .B(ram[3718]), .A(ram[3734]), .S(n12624), .Y(n10041) );
  MUX2X1 U11371 ( .B(n10040), .A(n10037), .S(n12588), .Y(n10051) );
  MUX2X1 U11372 ( .B(ram[3686]), .A(ram[3702]), .S(n12664), .Y(n10045) );
  MUX2X1 U11373 ( .B(ram[3654]), .A(ram[3670]), .S(n12680), .Y(n10044) );
  MUX2X1 U11374 ( .B(ram[3622]), .A(ram[3638]), .S(n12632), .Y(n10048) );
  MUX2X1 U11375 ( .B(ram[3590]), .A(ram[3606]), .S(n12637), .Y(n10047) );
  MUX2X1 U11376 ( .B(n10046), .A(n10043), .S(n12585), .Y(n10050) );
  MUX2X1 U11377 ( .B(n10049), .A(n10034), .S(n12567), .Y(n10084) );
  MUX2X1 U11378 ( .B(ram[3558]), .A(ram[3574]), .S(n12638), .Y(n10054) );
  MUX2X1 U11379 ( .B(ram[3526]), .A(ram[3542]), .S(n12642), .Y(n10053) );
  MUX2X1 U11380 ( .B(ram[3494]), .A(ram[3510]), .S(n12642), .Y(n10057) );
  MUX2X1 U11381 ( .B(ram[3462]), .A(ram[3478]), .S(n12621), .Y(n10056) );
  MUX2X1 U11382 ( .B(n10055), .A(n10052), .S(mem_access_addr[2]), .Y(n10066)
         );
  MUX2X1 U11383 ( .B(ram[3430]), .A(ram[3446]), .S(n12671), .Y(n10060) );
  MUX2X1 U11384 ( .B(ram[3398]), .A(ram[3414]), .S(n12665), .Y(n10059) );
  MUX2X1 U11385 ( .B(ram[3366]), .A(ram[3382]), .S(n12644), .Y(n10063) );
  MUX2X1 U11386 ( .B(ram[3334]), .A(ram[3350]), .S(n12681), .Y(n10062) );
  MUX2X1 U11387 ( .B(n10061), .A(n10058), .S(mem_access_addr[2]), .Y(n10065)
         );
  MUX2X1 U11388 ( .B(ram[3302]), .A(ram[3318]), .S(n12636), .Y(n10069) );
  MUX2X1 U11389 ( .B(ram[3270]), .A(ram[3286]), .S(n12629), .Y(n10068) );
  MUX2X1 U11390 ( .B(ram[3238]), .A(ram[3254]), .S(n12630), .Y(n10072) );
  MUX2X1 U11391 ( .B(ram[3206]), .A(ram[3222]), .S(n12643), .Y(n10071) );
  MUX2X1 U11392 ( .B(n10070), .A(n10067), .S(n12575), .Y(n10081) );
  MUX2X1 U11393 ( .B(ram[3174]), .A(ram[3190]), .S(n12627), .Y(n10075) );
  MUX2X1 U11394 ( .B(ram[3142]), .A(ram[3158]), .S(n12672), .Y(n10074) );
  MUX2X1 U11395 ( .B(ram[3110]), .A(ram[3126]), .S(n12644), .Y(n10078) );
  MUX2X1 U11396 ( .B(ram[3078]), .A(ram[3094]), .S(n12669), .Y(n10077) );
  MUX2X1 U11397 ( .B(n10076), .A(n10073), .S(mem_access_addr[2]), .Y(n10080)
         );
  MUX2X1 U11398 ( .B(n10079), .A(n10064), .S(n12564), .Y(n10083) );
  MUX2X1 U11399 ( .B(ram[3046]), .A(ram[3062]), .S(n12627), .Y(n10087) );
  MUX2X1 U11400 ( .B(ram[3014]), .A(ram[3030]), .S(n12634), .Y(n10086) );
  MUX2X1 U11401 ( .B(ram[2982]), .A(ram[2998]), .S(n12636), .Y(n10090) );
  MUX2X1 U11402 ( .B(ram[2950]), .A(ram[2966]), .S(n12645), .Y(n10089) );
  MUX2X1 U11403 ( .B(n10088), .A(n10085), .S(n12581), .Y(n10099) );
  MUX2X1 U11404 ( .B(ram[2918]), .A(ram[2934]), .S(n12681), .Y(n10093) );
  MUX2X1 U11405 ( .B(ram[2886]), .A(ram[2902]), .S(n12643), .Y(n10092) );
  MUX2X1 U11406 ( .B(ram[2854]), .A(ram[2870]), .S(n12637), .Y(n10096) );
  MUX2X1 U11407 ( .B(ram[2822]), .A(ram[2838]), .S(n12683), .Y(n10095) );
  MUX2X1 U11408 ( .B(n10094), .A(n10091), .S(n12576), .Y(n10098) );
  MUX2X1 U11409 ( .B(ram[2790]), .A(ram[2806]), .S(n12628), .Y(n10102) );
  MUX2X1 U11410 ( .B(ram[2758]), .A(ram[2774]), .S(n12621), .Y(n10101) );
  MUX2X1 U11411 ( .B(ram[2726]), .A(ram[2742]), .S(n12639), .Y(n10105) );
  MUX2X1 U11412 ( .B(ram[2694]), .A(ram[2710]), .S(n12638), .Y(n10104) );
  MUX2X1 U11413 ( .B(n10103), .A(n10100), .S(n12585), .Y(n10114) );
  MUX2X1 U11414 ( .B(ram[2662]), .A(ram[2678]), .S(n12653), .Y(n10108) );
  MUX2X1 U11415 ( .B(ram[2630]), .A(ram[2646]), .S(n12683), .Y(n10107) );
  MUX2X1 U11416 ( .B(ram[2598]), .A(ram[2614]), .S(n12672), .Y(n10111) );
  MUX2X1 U11417 ( .B(ram[2566]), .A(ram[2582]), .S(n12642), .Y(n10110) );
  MUX2X1 U11418 ( .B(n10109), .A(n10106), .S(n12576), .Y(n10113) );
  MUX2X1 U11419 ( .B(n10112), .A(n10097), .S(n12565), .Y(n10147) );
  MUX2X1 U11420 ( .B(ram[2534]), .A(ram[2550]), .S(n12622), .Y(n10117) );
  MUX2X1 U11421 ( .B(ram[2502]), .A(ram[2518]), .S(n12638), .Y(n10116) );
  MUX2X1 U11422 ( .B(ram[2470]), .A(ram[2486]), .S(n12648), .Y(n10120) );
  MUX2X1 U11423 ( .B(ram[2438]), .A(ram[2454]), .S(n12660), .Y(n10119) );
  MUX2X1 U11424 ( .B(n10118), .A(n10115), .S(n12577), .Y(n10129) );
  MUX2X1 U11425 ( .B(ram[2406]), .A(ram[2422]), .S(mem_access_addr[0]), .Y(
        n10123) );
  MUX2X1 U11426 ( .B(ram[2374]), .A(ram[2390]), .S(n12639), .Y(n10122) );
  MUX2X1 U11427 ( .B(ram[2342]), .A(ram[2358]), .S(n12622), .Y(n10126) );
  MUX2X1 U11428 ( .B(ram[2310]), .A(ram[2326]), .S(n12674), .Y(n10125) );
  MUX2X1 U11429 ( .B(n10124), .A(n10121), .S(n12587), .Y(n10128) );
  MUX2X1 U11430 ( .B(ram[2278]), .A(ram[2294]), .S(n12627), .Y(n10132) );
  MUX2X1 U11431 ( .B(ram[2246]), .A(ram[2262]), .S(n12641), .Y(n10131) );
  MUX2X1 U11432 ( .B(ram[2214]), .A(ram[2230]), .S(n12628), .Y(n10135) );
  MUX2X1 U11433 ( .B(ram[2182]), .A(ram[2198]), .S(n12650), .Y(n10134) );
  MUX2X1 U11434 ( .B(n10133), .A(n10130), .S(n12578), .Y(n10144) );
  MUX2X1 U11435 ( .B(ram[2150]), .A(ram[2166]), .S(n12633), .Y(n10138) );
  MUX2X1 U11436 ( .B(ram[2118]), .A(ram[2134]), .S(n12661), .Y(n10137) );
  MUX2X1 U11437 ( .B(ram[2086]), .A(ram[2102]), .S(n12659), .Y(n10141) );
  MUX2X1 U11438 ( .B(ram[2054]), .A(ram[2070]), .S(n12629), .Y(n10140) );
  MUX2X1 U11439 ( .B(n10139), .A(n10136), .S(n12580), .Y(n10143) );
  MUX2X1 U11440 ( .B(n10142), .A(n10127), .S(n12565), .Y(n10146) );
  MUX2X1 U11441 ( .B(n10145), .A(n10082), .S(mem_access_addr[6]), .Y(n10275)
         );
  MUX2X1 U11442 ( .B(ram[2022]), .A(ram[2038]), .S(n12632), .Y(n10150) );
  MUX2X1 U11443 ( .B(ram[1990]), .A(ram[2006]), .S(n12671), .Y(n10149) );
  MUX2X1 U11444 ( .B(ram[1958]), .A(ram[1974]), .S(n12628), .Y(n10153) );
  MUX2X1 U11445 ( .B(ram[1926]), .A(ram[1942]), .S(n12621), .Y(n10152) );
  MUX2X1 U11446 ( .B(n10151), .A(n10148), .S(n12586), .Y(n10162) );
  MUX2X1 U11447 ( .B(ram[1894]), .A(ram[1910]), .S(n12646), .Y(n10156) );
  MUX2X1 U11448 ( .B(ram[1862]), .A(ram[1878]), .S(n12637), .Y(n10155) );
  MUX2X1 U11449 ( .B(ram[1830]), .A(ram[1846]), .S(n12650), .Y(n10159) );
  MUX2X1 U11450 ( .B(ram[1798]), .A(ram[1814]), .S(n12683), .Y(n10158) );
  MUX2X1 U11451 ( .B(n10157), .A(n10154), .S(mem_access_addr[2]), .Y(n10161)
         );
  MUX2X1 U11452 ( .B(ram[1766]), .A(ram[1782]), .S(n12656), .Y(n10165) );
  MUX2X1 U11453 ( .B(ram[1734]), .A(ram[1750]), .S(n12653), .Y(n10164) );
  MUX2X1 U11454 ( .B(ram[1702]), .A(ram[1718]), .S(n12635), .Y(n10168) );
  MUX2X1 U11455 ( .B(ram[1670]), .A(ram[1686]), .S(n12676), .Y(n10167) );
  MUX2X1 U11456 ( .B(n10166), .A(n10163), .S(n12584), .Y(n10177) );
  MUX2X1 U11457 ( .B(ram[1638]), .A(ram[1654]), .S(n12637), .Y(n10171) );
  MUX2X1 U11458 ( .B(ram[1606]), .A(ram[1622]), .S(mem_access_addr[0]), .Y(
        n10170) );
  MUX2X1 U11459 ( .B(ram[1574]), .A(ram[1590]), .S(n12636), .Y(n10174) );
  MUX2X1 U11460 ( .B(ram[1542]), .A(ram[1558]), .S(n12624), .Y(n10173) );
  MUX2X1 U11461 ( .B(n10172), .A(n10169), .S(n12586), .Y(n10176) );
  MUX2X1 U11462 ( .B(n10175), .A(n10160), .S(n12567), .Y(n10210) );
  MUX2X1 U11463 ( .B(ram[1510]), .A(ram[1526]), .S(n12632), .Y(n10180) );
  MUX2X1 U11464 ( .B(ram[1478]), .A(ram[1494]), .S(n12653), .Y(n10179) );
  MUX2X1 U11465 ( .B(ram[1446]), .A(ram[1462]), .S(n12638), .Y(n10183) );
  MUX2X1 U11466 ( .B(ram[1414]), .A(ram[1430]), .S(mem_access_addr[0]), .Y(
        n10182) );
  MUX2X1 U11467 ( .B(n10181), .A(n10178), .S(n12582), .Y(n10192) );
  MUX2X1 U11468 ( .B(ram[1382]), .A(ram[1398]), .S(n12683), .Y(n10186) );
  MUX2X1 U11469 ( .B(ram[1350]), .A(ram[1366]), .S(n12644), .Y(n10185) );
  MUX2X1 U11470 ( .B(ram[1318]), .A(ram[1334]), .S(n12679), .Y(n10189) );
  MUX2X1 U11471 ( .B(ram[1286]), .A(ram[1302]), .S(n12643), .Y(n10188) );
  MUX2X1 U11472 ( .B(n10187), .A(n10184), .S(n12588), .Y(n10191) );
  MUX2X1 U11473 ( .B(ram[1254]), .A(ram[1270]), .S(n12631), .Y(n10195) );
  MUX2X1 U11474 ( .B(ram[1222]), .A(ram[1238]), .S(n12648), .Y(n10194) );
  MUX2X1 U11475 ( .B(ram[1190]), .A(ram[1206]), .S(n12652), .Y(n10198) );
  MUX2X1 U11476 ( .B(ram[1158]), .A(ram[1174]), .S(n12665), .Y(n10197) );
  MUX2X1 U11477 ( .B(n10196), .A(n10193), .S(n12588), .Y(n10207) );
  MUX2X1 U11478 ( .B(ram[1126]), .A(ram[1142]), .S(n12682), .Y(n10201) );
  MUX2X1 U11479 ( .B(ram[1094]), .A(ram[1110]), .S(n12635), .Y(n10200) );
  MUX2X1 U11480 ( .B(ram[1062]), .A(ram[1078]), .S(n12626), .Y(n10204) );
  MUX2X1 U11481 ( .B(ram[1030]), .A(ram[1046]), .S(n12635), .Y(n10203) );
  MUX2X1 U11482 ( .B(n10202), .A(n10199), .S(n12585), .Y(n10206) );
  MUX2X1 U11483 ( .B(n10205), .A(n10190), .S(n12566), .Y(n10209) );
  MUX2X1 U11484 ( .B(ram[998]), .A(ram[1014]), .S(n12636), .Y(n10213) );
  MUX2X1 U11485 ( .B(ram[966]), .A(ram[982]), .S(n12622), .Y(n10212) );
  MUX2X1 U11486 ( .B(ram[934]), .A(ram[950]), .S(n12668), .Y(n10216) );
  MUX2X1 U11487 ( .B(ram[902]), .A(ram[918]), .S(n12631), .Y(n10215) );
  MUX2X1 U11488 ( .B(n10214), .A(n10211), .S(n12581), .Y(n10225) );
  MUX2X1 U11489 ( .B(ram[870]), .A(ram[886]), .S(n12623), .Y(n10219) );
  MUX2X1 U11490 ( .B(ram[838]), .A(ram[854]), .S(n12682), .Y(n10218) );
  MUX2X1 U11491 ( .B(ram[806]), .A(ram[822]), .S(n12628), .Y(n10222) );
  MUX2X1 U11492 ( .B(ram[774]), .A(ram[790]), .S(n12635), .Y(n10221) );
  MUX2X1 U11493 ( .B(n10220), .A(n10217), .S(mem_access_addr[2]), .Y(n10224)
         );
  MUX2X1 U11494 ( .B(ram[742]), .A(ram[758]), .S(n12639), .Y(n10228) );
  MUX2X1 U11495 ( .B(ram[710]), .A(ram[726]), .S(n12670), .Y(n10227) );
  MUX2X1 U11496 ( .B(ram[678]), .A(ram[694]), .S(n12627), .Y(n10231) );
  MUX2X1 U11497 ( .B(ram[646]), .A(ram[662]), .S(n12640), .Y(n10230) );
  MUX2X1 U11498 ( .B(n10229), .A(n10226), .S(n12586), .Y(n10240) );
  MUX2X1 U11499 ( .B(ram[614]), .A(ram[630]), .S(n12642), .Y(n10234) );
  MUX2X1 U11500 ( .B(ram[582]), .A(ram[598]), .S(n12657), .Y(n10233) );
  MUX2X1 U11501 ( .B(ram[550]), .A(ram[566]), .S(n12683), .Y(n10237) );
  MUX2X1 U11502 ( .B(ram[518]), .A(ram[534]), .S(n12654), .Y(n10236) );
  MUX2X1 U11503 ( .B(n10235), .A(n10232), .S(n12588), .Y(n10239) );
  MUX2X1 U11504 ( .B(n10238), .A(n10223), .S(n12564), .Y(n10273) );
  MUX2X1 U11505 ( .B(ram[486]), .A(ram[502]), .S(n12664), .Y(n10243) );
  MUX2X1 U11506 ( .B(ram[454]), .A(ram[470]), .S(n12669), .Y(n10242) );
  MUX2X1 U11507 ( .B(ram[422]), .A(ram[438]), .S(n12638), .Y(n10246) );
  MUX2X1 U11508 ( .B(ram[390]), .A(ram[406]), .S(n12622), .Y(n10245) );
  MUX2X1 U11509 ( .B(n10244), .A(n10241), .S(mem_access_addr[2]), .Y(n10255)
         );
  MUX2X1 U11510 ( .B(ram[358]), .A(ram[374]), .S(n12663), .Y(n10249) );
  MUX2X1 U11511 ( .B(ram[326]), .A(ram[342]), .S(n12649), .Y(n10248) );
  MUX2X1 U11512 ( .B(ram[294]), .A(ram[310]), .S(n12665), .Y(n10252) );
  MUX2X1 U11513 ( .B(ram[262]), .A(ram[278]), .S(n12622), .Y(n10251) );
  MUX2X1 U11514 ( .B(n10250), .A(n10247), .S(n12588), .Y(n10254) );
  MUX2X1 U11515 ( .B(ram[230]), .A(ram[246]), .S(n12660), .Y(n10258) );
  MUX2X1 U11516 ( .B(ram[198]), .A(ram[214]), .S(n12658), .Y(n10257) );
  MUX2X1 U11517 ( .B(ram[166]), .A(ram[182]), .S(n12635), .Y(n10261) );
  MUX2X1 U11518 ( .B(ram[134]), .A(ram[150]), .S(n12651), .Y(n10260) );
  MUX2X1 U11519 ( .B(n10259), .A(n10256), .S(n12588), .Y(n10270) );
  MUX2X1 U11520 ( .B(ram[102]), .A(ram[118]), .S(n12675), .Y(n10264) );
  MUX2X1 U11521 ( .B(ram[70]), .A(ram[86]), .S(n12647), .Y(n10263) );
  MUX2X1 U11522 ( .B(ram[38]), .A(ram[54]), .S(n12648), .Y(n10267) );
  MUX2X1 U11523 ( .B(ram[6]), .A(ram[22]), .S(n12676), .Y(n10266) );
  MUX2X1 U11524 ( .B(n10265), .A(n10262), .S(n12580), .Y(n10269) );
  MUX2X1 U11525 ( .B(n10268), .A(n10253), .S(n12564), .Y(n10272) );
  MUX2X1 U11526 ( .B(n10271), .A(n10208), .S(mem_access_addr[6]), .Y(n10274)
         );
  MUX2X1 U11527 ( .B(ram[4071]), .A(ram[4087]), .S(n12675), .Y(n10278) );
  MUX2X1 U11528 ( .B(ram[4039]), .A(ram[4055]), .S(n12668), .Y(n10277) );
  MUX2X1 U11529 ( .B(ram[4007]), .A(ram[4023]), .S(n12631), .Y(n10281) );
  MUX2X1 U11530 ( .B(ram[3975]), .A(ram[3991]), .S(n12653), .Y(n10280) );
  MUX2X1 U11531 ( .B(n10279), .A(n10276), .S(n12577), .Y(n10290) );
  MUX2X1 U11532 ( .B(ram[3943]), .A(ram[3959]), .S(n12625), .Y(n10284) );
  MUX2X1 U11533 ( .B(ram[3911]), .A(ram[3927]), .S(n12646), .Y(n10283) );
  MUX2X1 U11534 ( .B(ram[3879]), .A(ram[3895]), .S(n12659), .Y(n10287) );
  MUX2X1 U11535 ( .B(ram[3847]), .A(ram[3863]), .S(n12655), .Y(n10286) );
  MUX2X1 U11536 ( .B(n10285), .A(n10282), .S(n12588), .Y(n10289) );
  MUX2X1 U11537 ( .B(ram[3815]), .A(ram[3831]), .S(n12680), .Y(n10293) );
  MUX2X1 U11538 ( .B(ram[3783]), .A(ram[3799]), .S(n12666), .Y(n10292) );
  MUX2X1 U11539 ( .B(ram[3751]), .A(ram[3767]), .S(n12674), .Y(n10296) );
  MUX2X1 U11540 ( .B(ram[3719]), .A(ram[3735]), .S(n12628), .Y(n10295) );
  MUX2X1 U11541 ( .B(n10294), .A(n10291), .S(n12583), .Y(n10305) );
  MUX2X1 U11542 ( .B(ram[3687]), .A(ram[3703]), .S(n12635), .Y(n10299) );
  MUX2X1 U11543 ( .B(ram[3655]), .A(ram[3671]), .S(n12671), .Y(n10298) );
  MUX2X1 U11544 ( .B(ram[3623]), .A(ram[3639]), .S(n12626), .Y(n10302) );
  MUX2X1 U11545 ( .B(ram[3591]), .A(ram[3607]), .S(n12659), .Y(n10301) );
  MUX2X1 U11546 ( .B(n10300), .A(n10297), .S(n12580), .Y(n10304) );
  MUX2X1 U11547 ( .B(n10303), .A(n10288), .S(n12567), .Y(n10338) );
  MUX2X1 U11548 ( .B(ram[3559]), .A(ram[3575]), .S(n12679), .Y(n10308) );
  MUX2X1 U11549 ( .B(ram[3527]), .A(ram[3543]), .S(n12682), .Y(n10307) );
  MUX2X1 U11550 ( .B(ram[3495]), .A(ram[3511]), .S(n12657), .Y(n10311) );
  MUX2X1 U11551 ( .B(ram[3463]), .A(ram[3479]), .S(n12625), .Y(n10310) );
  MUX2X1 U11552 ( .B(n10309), .A(n10306), .S(n12582), .Y(n10320) );
  MUX2X1 U11553 ( .B(ram[3431]), .A(ram[3447]), .S(n12668), .Y(n10314) );
  MUX2X1 U11554 ( .B(ram[3399]), .A(ram[3415]), .S(n12674), .Y(n10313) );
  MUX2X1 U11555 ( .B(ram[3367]), .A(ram[3383]), .S(n12628), .Y(n10317) );
  MUX2X1 U11556 ( .B(ram[3335]), .A(ram[3351]), .S(n12627), .Y(n10316) );
  MUX2X1 U11557 ( .B(n10315), .A(n10312), .S(n12578), .Y(n10319) );
  MUX2X1 U11558 ( .B(ram[3303]), .A(ram[3319]), .S(n12652), .Y(n10323) );
  MUX2X1 U11559 ( .B(ram[3271]), .A(ram[3287]), .S(n12621), .Y(n10322) );
  MUX2X1 U11560 ( .B(ram[3239]), .A(ram[3255]), .S(n12635), .Y(n10326) );
  MUX2X1 U11561 ( .B(ram[3207]), .A(ram[3223]), .S(mem_access_addr[0]), .Y(
        n10325) );
  MUX2X1 U11562 ( .B(n10324), .A(n10321), .S(n12578), .Y(n10335) );
  MUX2X1 U11563 ( .B(ram[3175]), .A(ram[3191]), .S(n12682), .Y(n10329) );
  MUX2X1 U11564 ( .B(ram[3143]), .A(ram[3159]), .S(n12680), .Y(n10328) );
  MUX2X1 U11565 ( .B(ram[3111]), .A(ram[3127]), .S(n12681), .Y(n10332) );
  MUX2X1 U11566 ( .B(ram[3079]), .A(ram[3095]), .S(n12634), .Y(n10331) );
  MUX2X1 U11567 ( .B(n10330), .A(n10327), .S(n12584), .Y(n10334) );
  MUX2X1 U11568 ( .B(n10333), .A(n10318), .S(n12565), .Y(n10337) );
  MUX2X1 U11569 ( .B(ram[3047]), .A(ram[3063]), .S(n12628), .Y(n10341) );
  MUX2X1 U11570 ( .B(ram[3015]), .A(ram[3031]), .S(n12629), .Y(n10340) );
  MUX2X1 U11571 ( .B(ram[2983]), .A(ram[2999]), .S(n12652), .Y(n10344) );
  MUX2X1 U11572 ( .B(ram[2951]), .A(ram[2967]), .S(n12633), .Y(n10343) );
  MUX2X1 U11573 ( .B(n10342), .A(n10339), .S(n12587), .Y(n10353) );
  MUX2X1 U11574 ( .B(ram[2919]), .A(ram[2935]), .S(n12628), .Y(n10347) );
  MUX2X1 U11575 ( .B(ram[2887]), .A(ram[2903]), .S(n12641), .Y(n10346) );
  MUX2X1 U11576 ( .B(ram[2855]), .A(ram[2871]), .S(n12682), .Y(n10350) );
  MUX2X1 U11577 ( .B(ram[2823]), .A(ram[2839]), .S(n12624), .Y(n10349) );
  MUX2X1 U11578 ( .B(n10348), .A(n10345), .S(n12586), .Y(n10352) );
  MUX2X1 U11579 ( .B(ram[2791]), .A(ram[2807]), .S(n12652), .Y(n10356) );
  MUX2X1 U11580 ( .B(ram[2759]), .A(ram[2775]), .S(n12637), .Y(n10355) );
  MUX2X1 U11581 ( .B(ram[2727]), .A(ram[2743]), .S(n12637), .Y(n10359) );
  MUX2X1 U11582 ( .B(ram[2695]), .A(ram[2711]), .S(n12636), .Y(n10358) );
  MUX2X1 U11583 ( .B(n10357), .A(n10354), .S(n12576), .Y(n10368) );
  MUX2X1 U11584 ( .B(ram[2663]), .A(ram[2679]), .S(n12630), .Y(n10362) );
  MUX2X1 U11585 ( .B(ram[2631]), .A(ram[2647]), .S(n12623), .Y(n10361) );
  MUX2X1 U11586 ( .B(ram[2599]), .A(ram[2615]), .S(n12638), .Y(n10365) );
  MUX2X1 U11587 ( .B(ram[2567]), .A(ram[2583]), .S(n12622), .Y(n10364) );
  MUX2X1 U11588 ( .B(n10363), .A(n10360), .S(n12579), .Y(n10367) );
  MUX2X1 U11589 ( .B(n10366), .A(n10351), .S(n12567), .Y(n10401) );
  MUX2X1 U11590 ( .B(ram[2535]), .A(ram[2551]), .S(n12646), .Y(n10371) );
  MUX2X1 U11591 ( .B(ram[2503]), .A(ram[2519]), .S(n12637), .Y(n10370) );
  MUX2X1 U11592 ( .B(ram[2471]), .A(ram[2487]), .S(n12622), .Y(n10374) );
  MUX2X1 U11593 ( .B(ram[2439]), .A(ram[2455]), .S(n12681), .Y(n10373) );
  MUX2X1 U11594 ( .B(n10372), .A(n10369), .S(n12587), .Y(n10383) );
  MUX2X1 U11595 ( .B(ram[2407]), .A(ram[2423]), .S(n12621), .Y(n10377) );
  MUX2X1 U11596 ( .B(ram[2375]), .A(ram[2391]), .S(n12670), .Y(n10376) );
  MUX2X1 U11597 ( .B(ram[2343]), .A(ram[2359]), .S(n12677), .Y(n10380) );
  MUX2X1 U11598 ( .B(ram[2311]), .A(ram[2327]), .S(n12682), .Y(n10379) );
  MUX2X1 U11599 ( .B(n10378), .A(n10375), .S(n12586), .Y(n10382) );
  MUX2X1 U11600 ( .B(ram[2279]), .A(ram[2295]), .S(n12621), .Y(n10386) );
  MUX2X1 U11601 ( .B(ram[2247]), .A(ram[2263]), .S(n12659), .Y(n10385) );
  MUX2X1 U11602 ( .B(ram[2215]), .A(ram[2231]), .S(n12667), .Y(n10389) );
  MUX2X1 U11603 ( .B(ram[2183]), .A(ram[2199]), .S(n12652), .Y(n10388) );
  MUX2X1 U11604 ( .B(n10387), .A(n10384), .S(n12584), .Y(n10398) );
  MUX2X1 U11605 ( .B(ram[2151]), .A(ram[2167]), .S(n12625), .Y(n10392) );
  MUX2X1 U11606 ( .B(ram[2119]), .A(ram[2135]), .S(n12663), .Y(n10391) );
  MUX2X1 U11607 ( .B(ram[2087]), .A(ram[2103]), .S(n12629), .Y(n10395) );
  MUX2X1 U11608 ( .B(ram[2055]), .A(ram[2071]), .S(n12637), .Y(n10394) );
  MUX2X1 U11609 ( .B(n10393), .A(n10390), .S(n12589), .Y(n10397) );
  MUX2X1 U11610 ( .B(n10396), .A(n10381), .S(n12566), .Y(n10400) );
  MUX2X1 U11611 ( .B(n10399), .A(n10336), .S(mem_access_addr[6]), .Y(n10529)
         );
  MUX2X1 U11612 ( .B(ram[2023]), .A(ram[2039]), .S(n12662), .Y(n10404) );
  MUX2X1 U11613 ( .B(ram[1991]), .A(ram[2007]), .S(n12665), .Y(n10403) );
  MUX2X1 U11614 ( .B(ram[1959]), .A(ram[1975]), .S(n12626), .Y(n10407) );
  MUX2X1 U11615 ( .B(ram[1927]), .A(ram[1943]), .S(n12630), .Y(n10406) );
  MUX2X1 U11616 ( .B(n10405), .A(n10402), .S(n12587), .Y(n10416) );
  MUX2X1 U11617 ( .B(ram[1895]), .A(ram[1911]), .S(n12661), .Y(n10410) );
  MUX2X1 U11618 ( .B(ram[1863]), .A(ram[1879]), .S(n12683), .Y(n10409) );
  MUX2X1 U11619 ( .B(ram[1831]), .A(ram[1847]), .S(n12624), .Y(n10413) );
  MUX2X1 U11620 ( .B(ram[1799]), .A(ram[1815]), .S(n12683), .Y(n10412) );
  MUX2X1 U11621 ( .B(n10411), .A(n10408), .S(n12584), .Y(n10415) );
  MUX2X1 U11622 ( .B(ram[1767]), .A(ram[1783]), .S(n12630), .Y(n10419) );
  MUX2X1 U11623 ( .B(ram[1735]), .A(ram[1751]), .S(n12655), .Y(n10418) );
  MUX2X1 U11624 ( .B(ram[1703]), .A(ram[1719]), .S(n12671), .Y(n10422) );
  MUX2X1 U11625 ( .B(ram[1671]), .A(ram[1687]), .S(n12645), .Y(n10421) );
  MUX2X1 U11626 ( .B(n10420), .A(n10417), .S(n12589), .Y(n10431) );
  MUX2X1 U11627 ( .B(ram[1639]), .A(ram[1655]), .S(n12625), .Y(n10425) );
  MUX2X1 U11628 ( .B(ram[1607]), .A(ram[1623]), .S(n12667), .Y(n10424) );
  MUX2X1 U11629 ( .B(ram[1575]), .A(ram[1591]), .S(n12647), .Y(n10428) );
  MUX2X1 U11630 ( .B(ram[1543]), .A(ram[1559]), .S(n12673), .Y(n10427) );
  MUX2X1 U11631 ( .B(n10426), .A(n10423), .S(n12589), .Y(n10430) );
  MUX2X1 U11632 ( .B(n10429), .A(n10414), .S(n12565), .Y(n10464) );
  MUX2X1 U11633 ( .B(ram[1511]), .A(ram[1527]), .S(n12660), .Y(n10434) );
  MUX2X1 U11634 ( .B(ram[1479]), .A(ram[1495]), .S(n12636), .Y(n10433) );
  MUX2X1 U11635 ( .B(ram[1447]), .A(ram[1463]), .S(n12633), .Y(n10437) );
  MUX2X1 U11636 ( .B(ram[1415]), .A(ram[1431]), .S(n12662), .Y(n10436) );
  MUX2X1 U11637 ( .B(n10435), .A(n10432), .S(n12586), .Y(n10446) );
  MUX2X1 U11638 ( .B(ram[1383]), .A(ram[1399]), .S(n12653), .Y(n10440) );
  MUX2X1 U11639 ( .B(ram[1351]), .A(ram[1367]), .S(n12628), .Y(n10439) );
  MUX2X1 U11640 ( .B(ram[1319]), .A(ram[1335]), .S(n12672), .Y(n10443) );
  MUX2X1 U11641 ( .B(ram[1287]), .A(ram[1303]), .S(n12654), .Y(n10442) );
  MUX2X1 U11642 ( .B(n10441), .A(n10438), .S(n12589), .Y(n10445) );
  MUX2X1 U11643 ( .B(ram[1255]), .A(ram[1271]), .S(n12663), .Y(n10449) );
  MUX2X1 U11644 ( .B(ram[1223]), .A(ram[1239]), .S(n12674), .Y(n10448) );
  MUX2X1 U11645 ( .B(ram[1191]), .A(ram[1207]), .S(n12658), .Y(n10452) );
  MUX2X1 U11646 ( .B(ram[1159]), .A(ram[1175]), .S(n12665), .Y(n10451) );
  MUX2X1 U11647 ( .B(n10450), .A(n10447), .S(n12586), .Y(n10461) );
  MUX2X1 U11648 ( .B(ram[1127]), .A(ram[1143]), .S(n12654), .Y(n10455) );
  MUX2X1 U11649 ( .B(ram[1095]), .A(ram[1111]), .S(n12634), .Y(n10454) );
  MUX2X1 U11650 ( .B(ram[1063]), .A(ram[1079]), .S(n12646), .Y(n10458) );
  MUX2X1 U11651 ( .B(ram[1031]), .A(ram[1047]), .S(n12650), .Y(n10457) );
  MUX2X1 U11652 ( .B(n10456), .A(n10453), .S(n12589), .Y(n10460) );
  MUX2X1 U11653 ( .B(n10459), .A(n10444), .S(n12564), .Y(n10463) );
  MUX2X1 U11654 ( .B(ram[999]), .A(ram[1015]), .S(n12679), .Y(n10467) );
  MUX2X1 U11655 ( .B(ram[967]), .A(ram[983]), .S(n12662), .Y(n10466) );
  MUX2X1 U11656 ( .B(ram[935]), .A(ram[951]), .S(n12677), .Y(n10470) );
  MUX2X1 U11657 ( .B(ram[903]), .A(ram[919]), .S(n12646), .Y(n10469) );
  MUX2X1 U11658 ( .B(n10468), .A(n10465), .S(n12575), .Y(n10479) );
  MUX2X1 U11659 ( .B(ram[871]), .A(ram[887]), .S(n12672), .Y(n10473) );
  MUX2X1 U11660 ( .B(ram[839]), .A(ram[855]), .S(n12644), .Y(n10472) );
  MUX2X1 U11661 ( .B(ram[807]), .A(ram[823]), .S(n12659), .Y(n10476) );
  MUX2X1 U11662 ( .B(ram[775]), .A(ram[791]), .S(n12643), .Y(n10475) );
  MUX2X1 U11663 ( .B(n10474), .A(n10471), .S(n12589), .Y(n10478) );
  MUX2X1 U11664 ( .B(ram[743]), .A(ram[759]), .S(n12672), .Y(n10482) );
  MUX2X1 U11665 ( .B(ram[711]), .A(ram[727]), .S(n12641), .Y(n10481) );
  MUX2X1 U11666 ( .B(ram[679]), .A(ram[695]), .S(n12665), .Y(n10485) );
  MUX2X1 U11667 ( .B(ram[647]), .A(ram[663]), .S(n12626), .Y(n10484) );
  MUX2X1 U11668 ( .B(n10483), .A(n10480), .S(n12575), .Y(n10494) );
  MUX2X1 U11669 ( .B(ram[615]), .A(ram[631]), .S(n12676), .Y(n10488) );
  MUX2X1 U11670 ( .B(ram[583]), .A(ram[599]), .S(n12623), .Y(n10487) );
  MUX2X1 U11671 ( .B(ram[551]), .A(ram[567]), .S(n12637), .Y(n10491) );
  MUX2X1 U11672 ( .B(ram[519]), .A(ram[535]), .S(n12625), .Y(n10490) );
  MUX2X1 U11673 ( .B(n10489), .A(n10486), .S(n12575), .Y(n10493) );
  MUX2X1 U11674 ( .B(n10492), .A(n10477), .S(n12567), .Y(n10527) );
  MUX2X1 U11675 ( .B(ram[487]), .A(ram[503]), .S(n12621), .Y(n10497) );
  MUX2X1 U11676 ( .B(ram[455]), .A(ram[471]), .S(n12629), .Y(n10496) );
  MUX2X1 U11677 ( .B(ram[423]), .A(ram[439]), .S(n12627), .Y(n10500) );
  MUX2X1 U11678 ( .B(ram[391]), .A(ram[407]), .S(n12660), .Y(n10499) );
  MUX2X1 U11679 ( .B(n10498), .A(n10495), .S(n12578), .Y(n10509) );
  MUX2X1 U11680 ( .B(ram[359]), .A(ram[375]), .S(n12683), .Y(n10503) );
  MUX2X1 U11681 ( .B(ram[327]), .A(ram[343]), .S(n12623), .Y(n10502) );
  MUX2X1 U11682 ( .B(ram[295]), .A(ram[311]), .S(n12624), .Y(n10506) );
  MUX2X1 U11683 ( .B(ram[263]), .A(ram[279]), .S(n12651), .Y(n10505) );
  MUX2X1 U11684 ( .B(n10504), .A(n10501), .S(n12586), .Y(n10508) );
  MUX2X1 U11685 ( .B(ram[231]), .A(ram[247]), .S(n12659), .Y(n10512) );
  MUX2X1 U11686 ( .B(ram[199]), .A(ram[215]), .S(n12673), .Y(n10511) );
  MUX2X1 U11687 ( .B(ram[167]), .A(ram[183]), .S(n12632), .Y(n10515) );
  MUX2X1 U11688 ( .B(ram[135]), .A(ram[151]), .S(n12649), .Y(n10514) );
  MUX2X1 U11689 ( .B(n10513), .A(n10510), .S(n12584), .Y(n10524) );
  MUX2X1 U11690 ( .B(ram[103]), .A(ram[119]), .S(n12678), .Y(n10518) );
  MUX2X1 U11691 ( .B(ram[71]), .A(ram[87]), .S(n12670), .Y(n10517) );
  MUX2X1 U11692 ( .B(ram[39]), .A(ram[55]), .S(n12651), .Y(n10521) );
  MUX2X1 U11693 ( .B(ram[7]), .A(ram[23]), .S(n12681), .Y(n10520) );
  MUX2X1 U11694 ( .B(n10519), .A(n10516), .S(n12586), .Y(n10523) );
  MUX2X1 U11695 ( .B(n10522), .A(n10507), .S(n12567), .Y(n10526) );
  MUX2X1 U11696 ( .B(n10525), .A(n10462), .S(mem_access_addr[6]), .Y(n10528)
         );
  MUX2X1 U11697 ( .B(ram[4072]), .A(ram[4088]), .S(n12625), .Y(n10532) );
  MUX2X1 U11698 ( .B(ram[4040]), .A(ram[4056]), .S(n12644), .Y(n10531) );
  MUX2X1 U11699 ( .B(ram[4008]), .A(ram[4024]), .S(n12622), .Y(n10535) );
  MUX2X1 U11700 ( .B(ram[3976]), .A(ram[3992]), .S(n12651), .Y(n10534) );
  MUX2X1 U11701 ( .B(n10533), .A(n10530), .S(n12577), .Y(n10544) );
  MUX2X1 U11702 ( .B(ram[3944]), .A(ram[3960]), .S(n12646), .Y(n10538) );
  MUX2X1 U11703 ( .B(ram[3912]), .A(ram[3928]), .S(n12631), .Y(n10537) );
  MUX2X1 U11704 ( .B(ram[3880]), .A(ram[3896]), .S(n12680), .Y(n10541) );
  MUX2X1 U11705 ( .B(ram[3848]), .A(ram[3864]), .S(n12647), .Y(n10540) );
  MUX2X1 U11706 ( .B(n10539), .A(n10536), .S(n12575), .Y(n10543) );
  MUX2X1 U11707 ( .B(ram[3816]), .A(ram[3832]), .S(n12630), .Y(n10547) );
  MUX2X1 U11708 ( .B(ram[3784]), .A(ram[3800]), .S(n12676), .Y(n10546) );
  MUX2X1 U11709 ( .B(ram[3752]), .A(ram[3768]), .S(n12629), .Y(n10550) );
  MUX2X1 U11710 ( .B(ram[3720]), .A(ram[3736]), .S(n12657), .Y(n10549) );
  MUX2X1 U11711 ( .B(n10548), .A(n10545), .S(n12587), .Y(n10559) );
  MUX2X1 U11712 ( .B(ram[3688]), .A(ram[3704]), .S(n12633), .Y(n10553) );
  MUX2X1 U11713 ( .B(ram[3656]), .A(ram[3672]), .S(n12621), .Y(n10552) );
  MUX2X1 U11714 ( .B(ram[3624]), .A(ram[3640]), .S(n12669), .Y(n10556) );
  MUX2X1 U11715 ( .B(ram[3592]), .A(ram[3608]), .S(n12623), .Y(n10555) );
  MUX2X1 U11716 ( .B(n10554), .A(n10551), .S(n12575), .Y(n10558) );
  MUX2X1 U11717 ( .B(n10557), .A(n10542), .S(n12567), .Y(n10592) );
  MUX2X1 U11718 ( .B(ram[3560]), .A(ram[3576]), .S(n12653), .Y(n10562) );
  MUX2X1 U11719 ( .B(ram[3528]), .A(ram[3544]), .S(n12674), .Y(n10561) );
  MUX2X1 U11720 ( .B(ram[3496]), .A(ram[3512]), .S(n12625), .Y(n10565) );
  MUX2X1 U11721 ( .B(ram[3464]), .A(ram[3480]), .S(n12630), .Y(n10564) );
  MUX2X1 U11722 ( .B(n10563), .A(n10560), .S(n12587), .Y(n10574) );
  MUX2X1 U11723 ( .B(ram[3432]), .A(ram[3448]), .S(n12654), .Y(n10568) );
  MUX2X1 U11724 ( .B(ram[3400]), .A(ram[3416]), .S(n12679), .Y(n10567) );
  MUX2X1 U11725 ( .B(ram[3368]), .A(ram[3384]), .S(n12627), .Y(n10571) );
  MUX2X1 U11726 ( .B(ram[3336]), .A(ram[3352]), .S(n12645), .Y(n10570) );
  MUX2X1 U11727 ( .B(n10569), .A(n10566), .S(mem_access_addr[2]), .Y(n10573)
         );
  MUX2X1 U11728 ( .B(ram[3304]), .A(ram[3320]), .S(n12653), .Y(n10577) );
  MUX2X1 U11729 ( .B(ram[3272]), .A(ram[3288]), .S(n12664), .Y(n10576) );
  MUX2X1 U11730 ( .B(ram[3240]), .A(ram[3256]), .S(n12631), .Y(n10580) );
  MUX2X1 U11731 ( .B(ram[3208]), .A(ram[3224]), .S(n12673), .Y(n10579) );
  MUX2X1 U11732 ( .B(n10578), .A(n10575), .S(n12583), .Y(n10589) );
  MUX2X1 U11733 ( .B(ram[3176]), .A(ram[3192]), .S(n12657), .Y(n10583) );
  MUX2X1 U11734 ( .B(ram[3144]), .A(ram[3160]), .S(n12632), .Y(n10582) );
  MUX2X1 U11735 ( .B(ram[3112]), .A(ram[3128]), .S(n12678), .Y(n10586) );
  MUX2X1 U11736 ( .B(ram[3080]), .A(ram[3096]), .S(n12651), .Y(n10585) );
  MUX2X1 U11737 ( .B(n10584), .A(n10581), .S(n12580), .Y(n10588) );
  MUX2X1 U11738 ( .B(n10587), .A(n10572), .S(n12566), .Y(n10591) );
  MUX2X1 U11739 ( .B(ram[3048]), .A(ram[3064]), .S(n12650), .Y(n10595) );
  MUX2X1 U11740 ( .B(ram[3016]), .A(ram[3032]), .S(n12678), .Y(n10594) );
  MUX2X1 U11741 ( .B(ram[2984]), .A(ram[3000]), .S(n12636), .Y(n10598) );
  MUX2X1 U11742 ( .B(ram[2952]), .A(ram[2968]), .S(n12649), .Y(n10597) );
  MUX2X1 U11743 ( .B(n10596), .A(n10593), .S(n12589), .Y(n10607) );
  MUX2X1 U11744 ( .B(ram[2920]), .A(ram[2936]), .S(n12656), .Y(n10601) );
  MUX2X1 U11745 ( .B(ram[2888]), .A(ram[2904]), .S(n12624), .Y(n10600) );
  MUX2X1 U11746 ( .B(ram[2856]), .A(ram[2872]), .S(n12622), .Y(n10604) );
  MUX2X1 U11747 ( .B(ram[2824]), .A(ram[2840]), .S(n12648), .Y(n10603) );
  MUX2X1 U11748 ( .B(n10602), .A(n10599), .S(n12581), .Y(n10606) );
  MUX2X1 U11749 ( .B(ram[2792]), .A(ram[2808]), .S(n12647), .Y(n10610) );
  MUX2X1 U11750 ( .B(ram[2760]), .A(ram[2776]), .S(n12649), .Y(n10609) );
  MUX2X1 U11751 ( .B(ram[2728]), .A(ram[2744]), .S(n12652), .Y(n10613) );
  MUX2X1 U11752 ( .B(ram[2696]), .A(ram[2712]), .S(n12638), .Y(n10612) );
  MUX2X1 U11753 ( .B(n10611), .A(n10608), .S(n12587), .Y(n10622) );
  MUX2X1 U11754 ( .B(ram[2664]), .A(ram[2680]), .S(n12663), .Y(n10616) );
  MUX2X1 U11755 ( .B(ram[2632]), .A(ram[2648]), .S(n12634), .Y(n10615) );
  MUX2X1 U11756 ( .B(ram[2600]), .A(ram[2616]), .S(n12654), .Y(n10619) );
  MUX2X1 U11757 ( .B(ram[2568]), .A(ram[2584]), .S(n12679), .Y(n10618) );
  MUX2X1 U11758 ( .B(n10617), .A(n10614), .S(n12585), .Y(n10621) );
  MUX2X1 U11759 ( .B(n10620), .A(n10605), .S(n12566), .Y(n10655) );
  MUX2X1 U11760 ( .B(ram[2536]), .A(ram[2552]), .S(n12626), .Y(n10625) );
  MUX2X1 U11761 ( .B(ram[2504]), .A(ram[2520]), .S(n12675), .Y(n10624) );
  MUX2X1 U11762 ( .B(ram[2472]), .A(ram[2488]), .S(n12626), .Y(n10628) );
  MUX2X1 U11763 ( .B(ram[2440]), .A(ram[2456]), .S(n12656), .Y(n10627) );
  MUX2X1 U11764 ( .B(n10626), .A(n10623), .S(n12587), .Y(n10637) );
  MUX2X1 U11765 ( .B(ram[2408]), .A(ram[2424]), .S(n12682), .Y(n10631) );
  MUX2X1 U11766 ( .B(ram[2376]), .A(ram[2392]), .S(n12651), .Y(n10630) );
  MUX2X1 U11767 ( .B(ram[2344]), .A(ram[2360]), .S(n12631), .Y(n10634) );
  MUX2X1 U11768 ( .B(ram[2312]), .A(ram[2328]), .S(n12683), .Y(n10633) );
  MUX2X1 U11769 ( .B(n10632), .A(n10629), .S(mem_access_addr[2]), .Y(n10636)
         );
  MUX2X1 U11770 ( .B(ram[2280]), .A(ram[2296]), .S(n12648), .Y(n10640) );
  MUX2X1 U11771 ( .B(ram[2248]), .A(ram[2264]), .S(n12633), .Y(n10639) );
  MUX2X1 U11772 ( .B(ram[2216]), .A(ram[2232]), .S(n12626), .Y(n10643) );
  MUX2X1 U11773 ( .B(ram[2184]), .A(ram[2200]), .S(n12635), .Y(n10642) );
  MUX2X1 U11774 ( .B(n10641), .A(n10638), .S(n12575), .Y(n10652) );
  MUX2X1 U11775 ( .B(ram[2152]), .A(ram[2168]), .S(n12660), .Y(n10646) );
  MUX2X1 U11776 ( .B(ram[2120]), .A(ram[2136]), .S(n12643), .Y(n10645) );
  MUX2X1 U11777 ( .B(ram[2088]), .A(ram[2104]), .S(n12623), .Y(n10649) );
  MUX2X1 U11778 ( .B(ram[2056]), .A(ram[2072]), .S(n12645), .Y(n10648) );
  MUX2X1 U11779 ( .B(n10647), .A(n10644), .S(n12578), .Y(n10651) );
  MUX2X1 U11780 ( .B(n10650), .A(n10635), .S(n12564), .Y(n10654) );
  MUX2X1 U11781 ( .B(n10653), .A(n10590), .S(mem_access_addr[6]), .Y(n10783)
         );
  MUX2X1 U11782 ( .B(ram[2024]), .A(ram[2040]), .S(n12637), .Y(n10658) );
  MUX2X1 U11783 ( .B(ram[1992]), .A(ram[2008]), .S(n12655), .Y(n10657) );
  MUX2X1 U11784 ( .B(ram[1960]), .A(ram[1976]), .S(n12666), .Y(n10661) );
  MUX2X1 U11785 ( .B(ram[1928]), .A(ram[1944]), .S(n12679), .Y(n10660) );
  MUX2X1 U11786 ( .B(n10659), .A(n10656), .S(n12589), .Y(n10670) );
  MUX2X1 U11787 ( .B(ram[1896]), .A(ram[1912]), .S(n12670), .Y(n10664) );
  MUX2X1 U11788 ( .B(ram[1864]), .A(ram[1880]), .S(n12624), .Y(n10663) );
  MUX2X1 U11789 ( .B(ram[1832]), .A(ram[1848]), .S(n12679), .Y(n10667) );
  MUX2X1 U11790 ( .B(ram[1800]), .A(ram[1816]), .S(n12681), .Y(n10666) );
  MUX2X1 U11791 ( .B(n10665), .A(n10662), .S(n12587), .Y(n10669) );
  MUX2X1 U11792 ( .B(ram[1768]), .A(ram[1784]), .S(n12668), .Y(n10673) );
  MUX2X1 U11793 ( .B(ram[1736]), .A(ram[1752]), .S(n12673), .Y(n10672) );
  MUX2X1 U11794 ( .B(ram[1704]), .A(ram[1720]), .S(n12652), .Y(n10676) );
  MUX2X1 U11795 ( .B(ram[1672]), .A(ram[1688]), .S(n12667), .Y(n10675) );
  MUX2X1 U11796 ( .B(n10674), .A(n10671), .S(n12589), .Y(n10685) );
  MUX2X1 U11797 ( .B(ram[1640]), .A(ram[1656]), .S(n12632), .Y(n10679) );
  MUX2X1 U11798 ( .B(ram[1608]), .A(ram[1624]), .S(n12644), .Y(n10678) );
  MUX2X1 U11799 ( .B(ram[1576]), .A(ram[1592]), .S(n12638), .Y(n10682) );
  MUX2X1 U11800 ( .B(ram[1544]), .A(ram[1560]), .S(n12668), .Y(n10681) );
  MUX2X1 U11801 ( .B(n10680), .A(n10677), .S(n12577), .Y(n10684) );
  MUX2X1 U11802 ( .B(n10683), .A(n10668), .S(n12565), .Y(n10718) );
  MUX2X1 U11803 ( .B(ram[1512]), .A(ram[1528]), .S(n12658), .Y(n10688) );
  MUX2X1 U11804 ( .B(ram[1480]), .A(ram[1496]), .S(n12621), .Y(n10687) );
  MUX2X1 U11805 ( .B(ram[1448]), .A(ram[1464]), .S(n12640), .Y(n10691) );
  MUX2X1 U11806 ( .B(ram[1416]), .A(ram[1432]), .S(n12664), .Y(n10690) );
  MUX2X1 U11807 ( .B(n10689), .A(n10686), .S(n12586), .Y(n10700) );
  MUX2X1 U11808 ( .B(ram[1384]), .A(ram[1400]), .S(n12645), .Y(n10694) );
  MUX2X1 U11809 ( .B(ram[1352]), .A(ram[1368]), .S(n12671), .Y(n10693) );
  MUX2X1 U11810 ( .B(ram[1320]), .A(ram[1336]), .S(n12666), .Y(n10697) );
  MUX2X1 U11811 ( .B(ram[1288]), .A(ram[1304]), .S(n12673), .Y(n10696) );
  MUX2X1 U11812 ( .B(n10695), .A(n10692), .S(n12588), .Y(n10699) );
  MUX2X1 U11813 ( .B(ram[1256]), .A(ram[1272]), .S(n12655), .Y(n10703) );
  MUX2X1 U11814 ( .B(ram[1224]), .A(ram[1240]), .S(n12656), .Y(n10702) );
  MUX2X1 U11815 ( .B(ram[1192]), .A(ram[1208]), .S(n12662), .Y(n10706) );
  MUX2X1 U11816 ( .B(ram[1160]), .A(ram[1176]), .S(n12673), .Y(n10705) );
  MUX2X1 U11817 ( .B(n10704), .A(n10701), .S(n12581), .Y(n10715) );
  MUX2X1 U11818 ( .B(ram[1128]), .A(ram[1144]), .S(n12660), .Y(n10709) );
  MUX2X1 U11819 ( .B(ram[1096]), .A(ram[1112]), .S(n12632), .Y(n10708) );
  MUX2X1 U11820 ( .B(ram[1064]), .A(ram[1080]), .S(n12656), .Y(n10712) );
  MUX2X1 U11821 ( .B(ram[1032]), .A(ram[1048]), .S(n12646), .Y(n10711) );
  MUX2X1 U11822 ( .B(n10710), .A(n10707), .S(n12584), .Y(n10714) );
  MUX2X1 U11823 ( .B(n10713), .A(n10698), .S(n12565), .Y(n10717) );
  MUX2X1 U11824 ( .B(ram[1000]), .A(ram[1016]), .S(n12668), .Y(n10721) );
  MUX2X1 U11825 ( .B(ram[968]), .A(ram[984]), .S(n12679), .Y(n10720) );
  MUX2X1 U11826 ( .B(ram[936]), .A(ram[952]), .S(n12677), .Y(n10724) );
  MUX2X1 U11827 ( .B(ram[904]), .A(ram[920]), .S(n12645), .Y(n10723) );
  MUX2X1 U11828 ( .B(n10722), .A(n10719), .S(n12582), .Y(n10733) );
  MUX2X1 U11829 ( .B(ram[872]), .A(ram[888]), .S(n12633), .Y(n10727) );
  MUX2X1 U11830 ( .B(ram[840]), .A(ram[856]), .S(n12635), .Y(n10726) );
  MUX2X1 U11831 ( .B(ram[808]), .A(ram[824]), .S(n12626), .Y(n10730) );
  MUX2X1 U11832 ( .B(ram[776]), .A(ram[792]), .S(n12683), .Y(n10729) );
  MUX2X1 U11833 ( .B(n10728), .A(n10725), .S(n12588), .Y(n10732) );
  MUX2X1 U11834 ( .B(ram[744]), .A(ram[760]), .S(n12634), .Y(n10736) );
  MUX2X1 U11835 ( .B(ram[712]), .A(ram[728]), .S(n12625), .Y(n10735) );
  MUX2X1 U11836 ( .B(ram[680]), .A(ram[696]), .S(n12631), .Y(n10739) );
  MUX2X1 U11837 ( .B(ram[648]), .A(ram[664]), .S(n12621), .Y(n10738) );
  MUX2X1 U11838 ( .B(n10737), .A(n10734), .S(n12585), .Y(n10748) );
  MUX2X1 U11839 ( .B(ram[616]), .A(ram[632]), .S(n12636), .Y(n10742) );
  MUX2X1 U11840 ( .B(ram[584]), .A(ram[600]), .S(n12626), .Y(n10741) );
  MUX2X1 U11841 ( .B(ram[552]), .A(ram[568]), .S(n12635), .Y(n10745) );
  MUX2X1 U11842 ( .B(ram[520]), .A(ram[536]), .S(n12683), .Y(n10744) );
  MUX2X1 U11843 ( .B(n10743), .A(n10740), .S(n12578), .Y(n10747) );
  MUX2X1 U11844 ( .B(n10746), .A(n10731), .S(n12566), .Y(n10781) );
  MUX2X1 U11845 ( .B(ram[488]), .A(ram[504]), .S(n12648), .Y(n10751) );
  MUX2X1 U11846 ( .B(ram[456]), .A(ram[472]), .S(n12665), .Y(n10750) );
  MUX2X1 U11847 ( .B(ram[424]), .A(ram[440]), .S(n12663), .Y(n10754) );
  MUX2X1 U11848 ( .B(ram[392]), .A(ram[408]), .S(n12658), .Y(n10753) );
  MUX2X1 U11849 ( .B(n10752), .A(n10749), .S(n12587), .Y(n10763) );
  MUX2X1 U11850 ( .B(ram[360]), .A(ram[376]), .S(n12680), .Y(n10757) );
  MUX2X1 U11851 ( .B(ram[328]), .A(ram[344]), .S(n12639), .Y(n10756) );
  MUX2X1 U11852 ( .B(ram[296]), .A(ram[312]), .S(n12640), .Y(n10760) );
  MUX2X1 U11853 ( .B(ram[264]), .A(ram[280]), .S(n12640), .Y(n10759) );
  MUX2X1 U11854 ( .B(n10758), .A(n10755), .S(n12585), .Y(n10762) );
  MUX2X1 U11855 ( .B(ram[232]), .A(ram[248]), .S(n12643), .Y(n10766) );
  MUX2X1 U11856 ( .B(ram[200]), .A(ram[216]), .S(n12651), .Y(n10765) );
  MUX2X1 U11857 ( .B(ram[168]), .A(ram[184]), .S(n12675), .Y(n10769) );
  MUX2X1 U11858 ( .B(ram[136]), .A(ram[152]), .S(n12665), .Y(n10768) );
  MUX2X1 U11859 ( .B(n10767), .A(n10764), .S(n12588), .Y(n10778) );
  MUX2X1 U11860 ( .B(ram[104]), .A(ram[120]), .S(n12677), .Y(n10772) );
  MUX2X1 U11861 ( .B(ram[72]), .A(ram[88]), .S(mem_access_addr[0]), .Y(n10771)
         );
  MUX2X1 U11862 ( .B(ram[40]), .A(ram[56]), .S(n12674), .Y(n10775) );
  MUX2X1 U11863 ( .B(ram[8]), .A(ram[24]), .S(n12623), .Y(n10774) );
  MUX2X1 U11864 ( .B(n10773), .A(n10770), .S(n12575), .Y(n10777) );
  MUX2X1 U11865 ( .B(n10776), .A(n10761), .S(n12564), .Y(n10780) );
  MUX2X1 U11866 ( .B(n10779), .A(n10716), .S(mem_access_addr[6]), .Y(n10782)
         );
  MUX2X1 U11867 ( .B(ram[4073]), .A(ram[4089]), .S(n12628), .Y(n10786) );
  MUX2X1 U11868 ( .B(ram[4041]), .A(ram[4057]), .S(n12634), .Y(n10785) );
  MUX2X1 U11869 ( .B(ram[4009]), .A(ram[4025]), .S(n12629), .Y(n10789) );
  MUX2X1 U11870 ( .B(ram[3977]), .A(ram[3993]), .S(n12626), .Y(n10788) );
  MUX2X1 U11871 ( .B(n10787), .A(n10784), .S(n12577), .Y(n10798) );
  MUX2X1 U11872 ( .B(ram[3945]), .A(ram[3961]), .S(n12645), .Y(n10792) );
  MUX2X1 U11873 ( .B(ram[3913]), .A(ram[3929]), .S(n12669), .Y(n10791) );
  MUX2X1 U11874 ( .B(ram[3881]), .A(ram[3897]), .S(n12629), .Y(n10795) );
  MUX2X1 U11875 ( .B(ram[3849]), .A(ram[3865]), .S(n12674), .Y(n10794) );
  MUX2X1 U11876 ( .B(n10793), .A(n10790), .S(n12575), .Y(n10797) );
  MUX2X1 U11877 ( .B(ram[3817]), .A(ram[3833]), .S(n12623), .Y(n10801) );
  MUX2X1 U11878 ( .B(ram[3785]), .A(ram[3801]), .S(n12624), .Y(n10800) );
  MUX2X1 U11879 ( .B(ram[3753]), .A(ram[3769]), .S(n12630), .Y(n10804) );
  MUX2X1 U11880 ( .B(ram[3721]), .A(ram[3737]), .S(n12627), .Y(n10803) );
  MUX2X1 U11881 ( .B(n10802), .A(n10799), .S(n12577), .Y(n10813) );
  MUX2X1 U11882 ( .B(ram[3689]), .A(ram[3705]), .S(n12621), .Y(n10807) );
  MUX2X1 U11883 ( .B(ram[3657]), .A(ram[3673]), .S(mem_access_addr[0]), .Y(
        n10806) );
  MUX2X1 U11884 ( .B(ram[3625]), .A(ram[3641]), .S(n12636), .Y(n10810) );
  MUX2X1 U11885 ( .B(ram[3593]), .A(ram[3609]), .S(n12631), .Y(n10809) );
  MUX2X1 U11886 ( .B(n10808), .A(n10805), .S(n12579), .Y(n10812) );
  MUX2X1 U11887 ( .B(n10811), .A(n10796), .S(n12567), .Y(n10846) );
  MUX2X1 U11888 ( .B(ram[3561]), .A(ram[3577]), .S(n12635), .Y(n10816) );
  MUX2X1 U11889 ( .B(ram[3529]), .A(ram[3545]), .S(n12624), .Y(n10815) );
  MUX2X1 U11890 ( .B(ram[3497]), .A(ram[3513]), .S(n12623), .Y(n10819) );
  MUX2X1 U11891 ( .B(ram[3465]), .A(ram[3481]), .S(n12673), .Y(n10818) );
  MUX2X1 U11892 ( .B(n10817), .A(n10814), .S(n12587), .Y(n10828) );
  MUX2X1 U11893 ( .B(ram[3433]), .A(ram[3449]), .S(n12624), .Y(n10822) );
  MUX2X1 U11894 ( .B(ram[3401]), .A(ram[3417]), .S(n12636), .Y(n10821) );
  MUX2X1 U11895 ( .B(ram[3369]), .A(ram[3385]), .S(n12631), .Y(n10825) );
  MUX2X1 U11896 ( .B(ram[3337]), .A(ram[3353]), .S(n12629), .Y(n10824) );
  MUX2X1 U11897 ( .B(n10823), .A(n10820), .S(n12586), .Y(n10827) );
  MUX2X1 U11898 ( .B(ram[3305]), .A(ram[3321]), .S(n12655), .Y(n10831) );
  MUX2X1 U11899 ( .B(ram[3273]), .A(ram[3289]), .S(n12662), .Y(n10830) );
  MUX2X1 U11900 ( .B(ram[3241]), .A(ram[3257]), .S(n12632), .Y(n10834) );
  MUX2X1 U11901 ( .B(ram[3209]), .A(ram[3225]), .S(n12666), .Y(n10833) );
  MUX2X1 U11902 ( .B(n10832), .A(n10829), .S(n12575), .Y(n10843) );
  MUX2X1 U11903 ( .B(ram[3177]), .A(ram[3193]), .S(n12670), .Y(n10837) );
  MUX2X1 U11904 ( .B(ram[3145]), .A(ram[3161]), .S(n12678), .Y(n10836) );
  MUX2X1 U11905 ( .B(ram[3113]), .A(ram[3129]), .S(mem_access_addr[0]), .Y(
        n10840) );
  MUX2X1 U11906 ( .B(ram[3081]), .A(ram[3097]), .S(n12658), .Y(n10839) );
  MUX2X1 U11907 ( .B(n10838), .A(n10835), .S(n12587), .Y(n10842) );
  MUX2X1 U11908 ( .B(n10841), .A(n10826), .S(n12567), .Y(n10845) );
  MUX2X1 U11909 ( .B(ram[3049]), .A(ram[3065]), .S(n12626), .Y(n10849) );
  MUX2X1 U11910 ( .B(ram[3017]), .A(ram[3033]), .S(n12664), .Y(n10848) );
  MUX2X1 U11911 ( .B(ram[2985]), .A(ram[3001]), .S(n12654), .Y(n10852) );
  MUX2X1 U11912 ( .B(ram[2953]), .A(ram[2969]), .S(n12639), .Y(n10851) );
  MUX2X1 U11913 ( .B(n10850), .A(n10847), .S(n12575), .Y(n10861) );
  MUX2X1 U11914 ( .B(ram[2921]), .A(ram[2937]), .S(n12666), .Y(n10855) );
  MUX2X1 U11915 ( .B(ram[2889]), .A(ram[2905]), .S(n12648), .Y(n10854) );
  MUX2X1 U11916 ( .B(ram[2857]), .A(ram[2873]), .S(n12630), .Y(n10858) );
  MUX2X1 U11917 ( .B(ram[2825]), .A(ram[2841]), .S(n12628), .Y(n10857) );
  MUX2X1 U11918 ( .B(n10856), .A(n10853), .S(n12575), .Y(n10860) );
  MUX2X1 U11919 ( .B(ram[2793]), .A(ram[2809]), .S(n12631), .Y(n10864) );
  MUX2X1 U11920 ( .B(ram[2761]), .A(ram[2777]), .S(n12640), .Y(n10863) );
  MUX2X1 U11921 ( .B(ram[2729]), .A(ram[2745]), .S(n12642), .Y(n10867) );
  MUX2X1 U11922 ( .B(ram[2697]), .A(ram[2713]), .S(n12672), .Y(n10866) );
  MUX2X1 U11923 ( .B(n10865), .A(n10862), .S(n12575), .Y(n10876) );
  MUX2X1 U11924 ( .B(ram[2665]), .A(ram[2681]), .S(n12655), .Y(n10870) );
  MUX2X1 U11925 ( .B(ram[2633]), .A(ram[2649]), .S(n12680), .Y(n10869) );
  MUX2X1 U11926 ( .B(ram[2601]), .A(ram[2617]), .S(n12638), .Y(n10873) );
  MUX2X1 U11927 ( .B(ram[2569]), .A(ram[2585]), .S(n12673), .Y(n10872) );
  MUX2X1 U11928 ( .B(n10871), .A(n10868), .S(n12575), .Y(n10875) );
  MUX2X1 U11929 ( .B(n10874), .A(n10859), .S(n12564), .Y(n10909) );
  MUX2X1 U11930 ( .B(ram[2537]), .A(ram[2553]), .S(n12668), .Y(n10879) );
  MUX2X1 U11931 ( .B(ram[2505]), .A(ram[2521]), .S(n12676), .Y(n10878) );
  MUX2X1 U11932 ( .B(ram[2473]), .A(ram[2489]), .S(n12650), .Y(n10882) );
  MUX2X1 U11933 ( .B(ram[2441]), .A(ram[2457]), .S(n12656), .Y(n10881) );
  MUX2X1 U11934 ( .B(n10880), .A(n10877), .S(n12575), .Y(n10891) );
  MUX2X1 U11935 ( .B(ram[2409]), .A(ram[2425]), .S(n12627), .Y(n10885) );
  MUX2X1 U11936 ( .B(ram[2377]), .A(ram[2393]), .S(n12653), .Y(n10884) );
  MUX2X1 U11937 ( .B(ram[2345]), .A(ram[2361]), .S(n12655), .Y(n10888) );
  MUX2X1 U11938 ( .B(ram[2313]), .A(ram[2329]), .S(n12671), .Y(n10887) );
  MUX2X1 U11939 ( .B(n10886), .A(n10883), .S(n12575), .Y(n10890) );
  MUX2X1 U11940 ( .B(ram[2281]), .A(ram[2297]), .S(n12645), .Y(n10894) );
  MUX2X1 U11941 ( .B(ram[2249]), .A(ram[2265]), .S(n12626), .Y(n10893) );
  MUX2X1 U11942 ( .B(ram[2217]), .A(ram[2233]), .S(n12654), .Y(n10897) );
  MUX2X1 U11943 ( .B(ram[2185]), .A(ram[2201]), .S(n12675), .Y(n10896) );
  MUX2X1 U11944 ( .B(n10895), .A(n10892), .S(n12575), .Y(n10906) );
  MUX2X1 U11945 ( .B(ram[2153]), .A(ram[2169]), .S(n12629), .Y(n10900) );
  MUX2X1 U11946 ( .B(ram[2121]), .A(ram[2137]), .S(n12654), .Y(n10899) );
  MUX2X1 U11947 ( .B(ram[2089]), .A(ram[2105]), .S(n12622), .Y(n10903) );
  MUX2X1 U11948 ( .B(ram[2057]), .A(ram[2073]), .S(n12640), .Y(n10902) );
  MUX2X1 U11949 ( .B(n10901), .A(n10898), .S(n12575), .Y(n10905) );
  MUX2X1 U11950 ( .B(n10904), .A(n10889), .S(n12565), .Y(n10908) );
  MUX2X1 U11951 ( .B(n10907), .A(n10844), .S(mem_access_addr[6]), .Y(n11037)
         );
  MUX2X1 U11952 ( .B(ram[2025]), .A(ram[2041]), .S(n12679), .Y(n10912) );
  MUX2X1 U11953 ( .B(ram[1993]), .A(ram[2009]), .S(n12660), .Y(n10911) );
  MUX2X1 U11954 ( .B(ram[1961]), .A(ram[1977]), .S(n12652), .Y(n10915) );
  MUX2X1 U11955 ( .B(ram[1929]), .A(ram[1945]), .S(n12655), .Y(n10914) );
  MUX2X1 U11956 ( .B(n10913), .A(n10910), .S(n12575), .Y(n10924) );
  MUX2X1 U11957 ( .B(ram[1897]), .A(ram[1913]), .S(n12657), .Y(n10918) );
  MUX2X1 U11958 ( .B(ram[1865]), .A(ram[1881]), .S(n12657), .Y(n10917) );
  MUX2X1 U11959 ( .B(ram[1833]), .A(ram[1849]), .S(n12678), .Y(n10921) );
  MUX2X1 U11960 ( .B(ram[1801]), .A(ram[1817]), .S(n12652), .Y(n10920) );
  MUX2X1 U11961 ( .B(n10919), .A(n10916), .S(n12575), .Y(n10923) );
  MUX2X1 U11962 ( .B(ram[1769]), .A(ram[1785]), .S(n12650), .Y(n10927) );
  MUX2X1 U11963 ( .B(ram[1737]), .A(ram[1753]), .S(n12635), .Y(n10926) );
  MUX2X1 U11964 ( .B(ram[1705]), .A(ram[1721]), .S(n12627), .Y(n10930) );
  MUX2X1 U11965 ( .B(ram[1673]), .A(ram[1689]), .S(n12657), .Y(n10929) );
  MUX2X1 U11966 ( .B(n10928), .A(n10925), .S(n12575), .Y(n10939) );
  MUX2X1 U11967 ( .B(ram[1641]), .A(ram[1657]), .S(n12630), .Y(n10933) );
  MUX2X1 U11968 ( .B(ram[1609]), .A(ram[1625]), .S(n12677), .Y(n10932) );
  MUX2X1 U11969 ( .B(ram[1577]), .A(ram[1593]), .S(n12648), .Y(n10936) );
  MUX2X1 U11970 ( .B(ram[1545]), .A(ram[1561]), .S(n12657), .Y(n10935) );
  MUX2X1 U11971 ( .B(n10934), .A(n10931), .S(n12575), .Y(n10938) );
  MUX2X1 U11972 ( .B(n10937), .A(n10922), .S(n12567), .Y(n10972) );
  MUX2X1 U11973 ( .B(ram[1513]), .A(ram[1529]), .S(n12669), .Y(n10942) );
  MUX2X1 U11974 ( .B(ram[1481]), .A(ram[1497]), .S(n12653), .Y(n10941) );
  MUX2X1 U11975 ( .B(ram[1449]), .A(ram[1465]), .S(n12636), .Y(n10945) );
  MUX2X1 U11976 ( .B(ram[1417]), .A(ram[1433]), .S(n12636), .Y(n10944) );
  MUX2X1 U11977 ( .B(n10943), .A(n10940), .S(n12588), .Y(n10954) );
  MUX2X1 U11978 ( .B(ram[1385]), .A(ram[1401]), .S(n12639), .Y(n10948) );
  MUX2X1 U11979 ( .B(ram[1353]), .A(ram[1369]), .S(n12661), .Y(n10947) );
  MUX2X1 U11980 ( .B(ram[1321]), .A(ram[1337]), .S(n12650), .Y(n10951) );
  MUX2X1 U11981 ( .B(ram[1289]), .A(ram[1305]), .S(n12640), .Y(n10950) );
  MUX2X1 U11982 ( .B(n10949), .A(n10946), .S(n12587), .Y(n10953) );
  MUX2X1 U11983 ( .B(ram[1257]), .A(ram[1273]), .S(n12658), .Y(n10957) );
  MUX2X1 U11984 ( .B(ram[1225]), .A(ram[1241]), .S(n12623), .Y(n10956) );
  MUX2X1 U11985 ( .B(ram[1193]), .A(ram[1209]), .S(n12677), .Y(n10960) );
  MUX2X1 U11986 ( .B(ram[1161]), .A(ram[1177]), .S(n12660), .Y(n10959) );
  MUX2X1 U11987 ( .B(n10958), .A(n10955), .S(n12581), .Y(n10969) );
  MUX2X1 U11988 ( .B(ram[1129]), .A(ram[1145]), .S(n12623), .Y(n10963) );
  MUX2X1 U11989 ( .B(ram[1097]), .A(ram[1113]), .S(n12683), .Y(n10962) );
  MUX2X1 U11990 ( .B(ram[1065]), .A(ram[1081]), .S(n12645), .Y(n10966) );
  MUX2X1 U11991 ( .B(ram[1033]), .A(ram[1049]), .S(n12661), .Y(n10965) );
  MUX2X1 U11992 ( .B(n10964), .A(n10961), .S(n12587), .Y(n10968) );
  MUX2X1 U11993 ( .B(n10967), .A(n10952), .S(n12566), .Y(n10971) );
  MUX2X1 U11994 ( .B(ram[1001]), .A(ram[1017]), .S(n12679), .Y(n10975) );
  MUX2X1 U11995 ( .B(ram[969]), .A(ram[985]), .S(n12675), .Y(n10974) );
  MUX2X1 U11996 ( .B(ram[937]), .A(ram[953]), .S(n12680), .Y(n10978) );
  MUX2X1 U11997 ( .B(ram[905]), .A(ram[921]), .S(n12625), .Y(n10977) );
  MUX2X1 U11998 ( .B(n10976), .A(n10973), .S(n12576), .Y(n10987) );
  MUX2X1 U11999 ( .B(ram[873]), .A(ram[889]), .S(n12657), .Y(n10981) );
  MUX2X1 U12000 ( .B(ram[841]), .A(ram[857]), .S(n12625), .Y(n10980) );
  MUX2X1 U12001 ( .B(ram[809]), .A(ram[825]), .S(n12673), .Y(n10984) );
  MUX2X1 U12002 ( .B(ram[777]), .A(ram[793]), .S(n12647), .Y(n10983) );
  MUX2X1 U12003 ( .B(n10982), .A(n10979), .S(n12589), .Y(n10986) );
  MUX2X1 U12004 ( .B(ram[745]), .A(ram[761]), .S(n12623), .Y(n10990) );
  MUX2X1 U12005 ( .B(ram[713]), .A(ram[729]), .S(n12622), .Y(n10989) );
  MUX2X1 U12006 ( .B(ram[681]), .A(ram[697]), .S(n12638), .Y(n10993) );
  MUX2X1 U12007 ( .B(ram[649]), .A(ram[665]), .S(n12632), .Y(n10992) );
  MUX2X1 U12008 ( .B(n10991), .A(n10988), .S(n12578), .Y(n11002) );
  MUX2X1 U12009 ( .B(ram[617]), .A(ram[633]), .S(n12623), .Y(n10996) );
  MUX2X1 U12010 ( .B(ram[585]), .A(ram[601]), .S(n12645), .Y(n10995) );
  MUX2X1 U12011 ( .B(ram[553]), .A(ram[569]), .S(n12621), .Y(n10999) );
  MUX2X1 U12012 ( .B(ram[521]), .A(ram[537]), .S(n12660), .Y(n10998) );
  MUX2X1 U12013 ( .B(n10997), .A(n10994), .S(n12584), .Y(n11001) );
  MUX2X1 U12014 ( .B(n11000), .A(n10985), .S(n12567), .Y(n11035) );
  MUX2X1 U12015 ( .B(ram[489]), .A(ram[505]), .S(n12623), .Y(n11005) );
  MUX2X1 U12016 ( .B(ram[457]), .A(ram[473]), .S(n12644), .Y(n11004) );
  MUX2X1 U12017 ( .B(ram[425]), .A(ram[441]), .S(n12626), .Y(n11008) );
  MUX2X1 U12018 ( .B(ram[393]), .A(ram[409]), .S(n12649), .Y(n11007) );
  MUX2X1 U12019 ( .B(n11006), .A(n11003), .S(n12587), .Y(n11017) );
  MUX2X1 U12020 ( .B(ram[361]), .A(ram[377]), .S(n12645), .Y(n11011) );
  MUX2X1 U12021 ( .B(ram[329]), .A(ram[345]), .S(n12628), .Y(n11010) );
  MUX2X1 U12022 ( .B(ram[297]), .A(ram[313]), .S(n12635), .Y(n11014) );
  MUX2X1 U12023 ( .B(ram[265]), .A(ram[281]), .S(n12640), .Y(n11013) );
  MUX2X1 U12024 ( .B(n11012), .A(n11009), .S(n12585), .Y(n11016) );
  MUX2X1 U12025 ( .B(ram[233]), .A(ram[249]), .S(n12655), .Y(n11020) );
  MUX2X1 U12026 ( .B(ram[201]), .A(ram[217]), .S(n12665), .Y(n11019) );
  MUX2X1 U12027 ( .B(ram[169]), .A(ram[185]), .S(n12681), .Y(n11023) );
  MUX2X1 U12028 ( .B(ram[137]), .A(ram[153]), .S(n12648), .Y(n11022) );
  MUX2X1 U12029 ( .B(n11021), .A(n11018), .S(n12589), .Y(n11032) );
  MUX2X1 U12030 ( .B(ram[105]), .A(ram[121]), .S(n12671), .Y(n11026) );
  MUX2X1 U12031 ( .B(ram[73]), .A(ram[89]), .S(n12624), .Y(n11025) );
  MUX2X1 U12032 ( .B(ram[41]), .A(ram[57]), .S(n12679), .Y(n11029) );
  MUX2X1 U12033 ( .B(ram[9]), .A(ram[25]), .S(n12642), .Y(n11028) );
  MUX2X1 U12034 ( .B(n11027), .A(n11024), .S(n12576), .Y(n11031) );
  MUX2X1 U12035 ( .B(n11030), .A(n11015), .S(n12564), .Y(n11034) );
  MUX2X1 U12036 ( .B(n11033), .A(n10970), .S(mem_access_addr[6]), .Y(n11036)
         );
  MUX2X1 U12037 ( .B(ram[4074]), .A(ram[4090]), .S(n12626), .Y(n11040) );
  MUX2X1 U12038 ( .B(ram[4042]), .A(ram[4058]), .S(n12664), .Y(n11039) );
  MUX2X1 U12039 ( .B(ram[4010]), .A(ram[4026]), .S(n12635), .Y(n11043) );
  MUX2X1 U12040 ( .B(ram[3978]), .A(ram[3994]), .S(n12652), .Y(n11042) );
  MUX2X1 U12041 ( .B(n11041), .A(n11038), .S(n12578), .Y(n11052) );
  MUX2X1 U12042 ( .B(ram[3946]), .A(ram[3962]), .S(n12666), .Y(n11046) );
  MUX2X1 U12043 ( .B(ram[3914]), .A(ram[3930]), .S(n12667), .Y(n11045) );
  MUX2X1 U12044 ( .B(ram[3882]), .A(ram[3898]), .S(n12639), .Y(n11049) );
  MUX2X1 U12045 ( .B(ram[3850]), .A(ram[3866]), .S(n12651), .Y(n11048) );
  MUX2X1 U12046 ( .B(n11047), .A(n11044), .S(n12581), .Y(n11051) );
  MUX2X1 U12047 ( .B(ram[3818]), .A(ram[3834]), .S(n12650), .Y(n11055) );
  MUX2X1 U12048 ( .B(ram[3786]), .A(ram[3802]), .S(n12640), .Y(n11054) );
  MUX2X1 U12049 ( .B(ram[3754]), .A(ram[3770]), .S(n12634), .Y(n11058) );
  MUX2X1 U12050 ( .B(ram[3722]), .A(ram[3738]), .S(n12626), .Y(n11057) );
  MUX2X1 U12051 ( .B(n11056), .A(n11053), .S(n12576), .Y(n11067) );
  MUX2X1 U12052 ( .B(ram[3690]), .A(ram[3706]), .S(n12672), .Y(n11061) );
  MUX2X1 U12053 ( .B(ram[3658]), .A(ram[3674]), .S(n12631), .Y(n11060) );
  MUX2X1 U12054 ( .B(ram[3626]), .A(ram[3642]), .S(n12634), .Y(n11064) );
  MUX2X1 U12055 ( .B(ram[3594]), .A(ram[3610]), .S(n12632), .Y(n11063) );
  MUX2X1 U12056 ( .B(n11062), .A(n11059), .S(n12582), .Y(n11066) );
  MUX2X1 U12057 ( .B(n11065), .A(n11050), .S(n12564), .Y(n11100) );
  MUX2X1 U12058 ( .B(ram[3562]), .A(ram[3578]), .S(n12639), .Y(n11070) );
  MUX2X1 U12059 ( .B(ram[3530]), .A(ram[3546]), .S(n12672), .Y(n11069) );
  MUX2X1 U12060 ( .B(ram[3498]), .A(ram[3514]), .S(n12656), .Y(n11073) );
  MUX2X1 U12061 ( .B(ram[3466]), .A(ram[3482]), .S(n12675), .Y(n11072) );
  MUX2X1 U12062 ( .B(n11071), .A(n11068), .S(n12576), .Y(n11082) );
  MUX2X1 U12063 ( .B(ram[3434]), .A(ram[3450]), .S(mem_access_addr[0]), .Y(
        n11076) );
  MUX2X1 U12064 ( .B(ram[3402]), .A(ram[3418]), .S(n12655), .Y(n11075) );
  MUX2X1 U12065 ( .B(ram[3370]), .A(ram[3386]), .S(n12646), .Y(n11079) );
  MUX2X1 U12066 ( .B(ram[3338]), .A(ram[3354]), .S(n12681), .Y(n11078) );
  MUX2X1 U12067 ( .B(n11077), .A(n11074), .S(n12583), .Y(n11081) );
  MUX2X1 U12068 ( .B(ram[3306]), .A(ram[3322]), .S(n12669), .Y(n11085) );
  MUX2X1 U12069 ( .B(ram[3274]), .A(ram[3290]), .S(n12665), .Y(n11084) );
  MUX2X1 U12070 ( .B(ram[3242]), .A(ram[3258]), .S(n12625), .Y(n11088) );
  MUX2X1 U12071 ( .B(ram[3210]), .A(ram[3226]), .S(n12641), .Y(n11087) );
  MUX2X1 U12072 ( .B(n11086), .A(n11083), .S(n12584), .Y(n11097) );
  MUX2X1 U12073 ( .B(ram[3178]), .A(ram[3194]), .S(n12622), .Y(n11091) );
  MUX2X1 U12074 ( .B(ram[3146]), .A(ram[3162]), .S(n12640), .Y(n11090) );
  MUX2X1 U12075 ( .B(ram[3114]), .A(ram[3130]), .S(n12629), .Y(n11094) );
  MUX2X1 U12076 ( .B(ram[3082]), .A(ram[3098]), .S(n12675), .Y(n11093) );
  MUX2X1 U12077 ( .B(n11092), .A(n11089), .S(n12579), .Y(n11096) );
  MUX2X1 U12078 ( .B(n11095), .A(n11080), .S(n12565), .Y(n11099) );
  MUX2X1 U12079 ( .B(ram[3050]), .A(ram[3066]), .S(n12632), .Y(n11103) );
  MUX2X1 U12080 ( .B(ram[3018]), .A(ram[3034]), .S(n12653), .Y(n11102) );
  MUX2X1 U12081 ( .B(ram[2986]), .A(ram[3002]), .S(n12633), .Y(n11106) );
  MUX2X1 U12082 ( .B(ram[2954]), .A(ram[2970]), .S(n12646), .Y(n11105) );
  MUX2X1 U12083 ( .B(n11104), .A(n11101), .S(n12581), .Y(n11115) );
  MUX2X1 U12084 ( .B(ram[2922]), .A(ram[2938]), .S(n12627), .Y(n11109) );
  MUX2X1 U12085 ( .B(ram[2890]), .A(ram[2906]), .S(n12660), .Y(n11108) );
  MUX2X1 U12086 ( .B(ram[2858]), .A(ram[2874]), .S(n12644), .Y(n11112) );
  MUX2X1 U12087 ( .B(ram[2826]), .A(ram[2842]), .S(n12626), .Y(n11111) );
  MUX2X1 U12088 ( .B(n11110), .A(n11107), .S(n12577), .Y(n11114) );
  MUX2X1 U12089 ( .B(ram[2794]), .A(ram[2810]), .S(n12630), .Y(n11118) );
  MUX2X1 U12090 ( .B(ram[2762]), .A(ram[2778]), .S(n12629), .Y(n11117) );
  MUX2X1 U12091 ( .B(ram[2730]), .A(ram[2746]), .S(n12634), .Y(n11121) );
  MUX2X1 U12092 ( .B(ram[2698]), .A(ram[2714]), .S(n12637), .Y(n11120) );
  MUX2X1 U12093 ( .B(n11119), .A(n11116), .S(n12576), .Y(n11130) );
  MUX2X1 U12094 ( .B(ram[2666]), .A(ram[2682]), .S(n12650), .Y(n11124) );
  MUX2X1 U12095 ( .B(ram[2634]), .A(ram[2650]), .S(n12635), .Y(n11123) );
  MUX2X1 U12096 ( .B(ram[2602]), .A(ram[2618]), .S(n12633), .Y(n11127) );
  MUX2X1 U12097 ( .B(ram[2570]), .A(ram[2586]), .S(n12649), .Y(n11126) );
  MUX2X1 U12098 ( .B(n11125), .A(n11122), .S(n12585), .Y(n11129) );
  MUX2X1 U12099 ( .B(n11128), .A(n11113), .S(n12564), .Y(n11163) );
  MUX2X1 U12100 ( .B(ram[2538]), .A(ram[2554]), .S(n12674), .Y(n11133) );
  MUX2X1 U12101 ( .B(ram[2506]), .A(ram[2522]), .S(mem_access_addr[0]), .Y(
        n11132) );
  MUX2X1 U12102 ( .B(ram[2474]), .A(ram[2490]), .S(n12633), .Y(n11136) );
  MUX2X1 U12103 ( .B(ram[2442]), .A(ram[2458]), .S(n12637), .Y(n11135) );
  MUX2X1 U12104 ( .B(n11134), .A(n11131), .S(n12576), .Y(n11145) );
  MUX2X1 U12105 ( .B(ram[2410]), .A(ram[2426]), .S(n12672), .Y(n11139) );
  MUX2X1 U12106 ( .B(ram[2378]), .A(ram[2394]), .S(n12642), .Y(n11138) );
  MUX2X1 U12107 ( .B(ram[2346]), .A(ram[2362]), .S(n12637), .Y(n11142) );
  MUX2X1 U12108 ( .B(ram[2314]), .A(ram[2330]), .S(n12664), .Y(n11141) );
  MUX2X1 U12109 ( .B(n11140), .A(n11137), .S(n12588), .Y(n11144) );
  MUX2X1 U12110 ( .B(ram[2282]), .A(ram[2298]), .S(n12638), .Y(n11148) );
  MUX2X1 U12111 ( .B(ram[2250]), .A(ram[2266]), .S(n12621), .Y(n11147) );
  MUX2X1 U12112 ( .B(ram[2218]), .A(ram[2234]), .S(n12635), .Y(n11151) );
  MUX2X1 U12113 ( .B(ram[2186]), .A(ram[2202]), .S(n12625), .Y(n11150) );
  MUX2X1 U12114 ( .B(n11149), .A(n11146), .S(n12588), .Y(n11160) );
  MUX2X1 U12115 ( .B(ram[2154]), .A(ram[2170]), .S(n12658), .Y(n11154) );
  MUX2X1 U12116 ( .B(ram[2122]), .A(ram[2138]), .S(n12665), .Y(n11153) );
  MUX2X1 U12117 ( .B(ram[2090]), .A(ram[2106]), .S(n12655), .Y(n11157) );
  MUX2X1 U12118 ( .B(ram[2058]), .A(ram[2074]), .S(n12651), .Y(n11156) );
  MUX2X1 U12119 ( .B(n11155), .A(n11152), .S(n12578), .Y(n11159) );
  MUX2X1 U12120 ( .B(n11158), .A(n11143), .S(n12566), .Y(n11162) );
  MUX2X1 U12121 ( .B(n11161), .A(n11098), .S(mem_access_addr[6]), .Y(n11291)
         );
  MUX2X1 U12122 ( .B(ram[2026]), .A(ram[2042]), .S(n12671), .Y(n11166) );
  MUX2X1 U12123 ( .B(ram[1994]), .A(ram[2010]), .S(n12680), .Y(n11165) );
  MUX2X1 U12124 ( .B(ram[1962]), .A(ram[1978]), .S(n12624), .Y(n11169) );
  MUX2X1 U12125 ( .B(ram[1930]), .A(ram[1946]), .S(n12657), .Y(n11168) );
  MUX2X1 U12126 ( .B(n11167), .A(n11164), .S(n12582), .Y(n11178) );
  MUX2X1 U12127 ( .B(ram[1898]), .A(ram[1914]), .S(n12674), .Y(n11172) );
  MUX2X1 U12128 ( .B(ram[1866]), .A(ram[1882]), .S(n12642), .Y(n11171) );
  MUX2X1 U12129 ( .B(ram[1834]), .A(ram[1850]), .S(n12636), .Y(n11175) );
  MUX2X1 U12130 ( .B(ram[1802]), .A(ram[1818]), .S(n12643), .Y(n11174) );
  MUX2X1 U12131 ( .B(n11173), .A(n11170), .S(n12587), .Y(n11177) );
  MUX2X1 U12132 ( .B(ram[1770]), .A(ram[1786]), .S(n12652), .Y(n11181) );
  MUX2X1 U12133 ( .B(ram[1738]), .A(ram[1754]), .S(n12665), .Y(n11180) );
  MUX2X1 U12134 ( .B(ram[1706]), .A(ram[1722]), .S(n12626), .Y(n11184) );
  MUX2X1 U12135 ( .B(ram[1674]), .A(ram[1690]), .S(n12624), .Y(n11183) );
  MUX2X1 U12136 ( .B(n11182), .A(n11179), .S(n12577), .Y(n11193) );
  MUX2X1 U12137 ( .B(ram[1642]), .A(ram[1658]), .S(n12678), .Y(n11187) );
  MUX2X1 U12138 ( .B(ram[1610]), .A(ram[1626]), .S(n12677), .Y(n11186) );
  MUX2X1 U12139 ( .B(ram[1578]), .A(ram[1594]), .S(n12667), .Y(n11190) );
  MUX2X1 U12140 ( .B(ram[1546]), .A(ram[1562]), .S(n12666), .Y(n11189) );
  MUX2X1 U12141 ( .B(n11188), .A(n11185), .S(n12579), .Y(n11192) );
  MUX2X1 U12142 ( .B(n11191), .A(n11176), .S(n12564), .Y(n11226) );
  MUX2X1 U12143 ( .B(ram[1514]), .A(ram[1530]), .S(n12659), .Y(n11196) );
  MUX2X1 U12144 ( .B(ram[1482]), .A(ram[1498]), .S(n12668), .Y(n11195) );
  MUX2X1 U12145 ( .B(ram[1450]), .A(ram[1466]), .S(n12681), .Y(n11199) );
  MUX2X1 U12146 ( .B(ram[1418]), .A(ram[1434]), .S(n12673), .Y(n11198) );
  MUX2X1 U12147 ( .B(n11197), .A(n11194), .S(n12580), .Y(n11208) );
  MUX2X1 U12148 ( .B(ram[1386]), .A(ram[1402]), .S(n12634), .Y(n11202) );
  MUX2X1 U12149 ( .B(ram[1354]), .A(ram[1370]), .S(n12651), .Y(n11201) );
  MUX2X1 U12150 ( .B(ram[1322]), .A(ram[1338]), .S(n12646), .Y(n11205) );
  MUX2X1 U12151 ( .B(ram[1290]), .A(ram[1306]), .S(n12652), .Y(n11204) );
  MUX2X1 U12152 ( .B(n11203), .A(n11200), .S(n12583), .Y(n11207) );
  MUX2X1 U12153 ( .B(ram[1258]), .A(ram[1274]), .S(n12650), .Y(n11211) );
  MUX2X1 U12154 ( .B(ram[1226]), .A(ram[1242]), .S(n12630), .Y(n11210) );
  MUX2X1 U12155 ( .B(ram[1194]), .A(ram[1210]), .S(n12637), .Y(n11214) );
  MUX2X1 U12156 ( .B(ram[1162]), .A(ram[1178]), .S(n12629), .Y(n11213) );
  MUX2X1 U12157 ( .B(n11212), .A(n11209), .S(n12583), .Y(n11223) );
  MUX2X1 U12158 ( .B(ram[1130]), .A(ram[1146]), .S(n12627), .Y(n11217) );
  MUX2X1 U12159 ( .B(ram[1098]), .A(ram[1114]), .S(n12682), .Y(n11216) );
  MUX2X1 U12160 ( .B(ram[1066]), .A(ram[1082]), .S(n12653), .Y(n11220) );
  MUX2X1 U12161 ( .B(ram[1034]), .A(ram[1050]), .S(n12645), .Y(n11219) );
  MUX2X1 U12162 ( .B(n11218), .A(n11215), .S(n12584), .Y(n11222) );
  MUX2X1 U12163 ( .B(n11221), .A(n11206), .S(n12566), .Y(n11225) );
  MUX2X1 U12164 ( .B(ram[1002]), .A(ram[1018]), .S(n12634), .Y(n11229) );
  MUX2X1 U12165 ( .B(ram[970]), .A(ram[986]), .S(n12676), .Y(n11228) );
  MUX2X1 U12166 ( .B(ram[938]), .A(ram[954]), .S(n12635), .Y(n11232) );
  MUX2X1 U12167 ( .B(ram[906]), .A(ram[922]), .S(mem_access_addr[0]), .Y(
        n11231) );
  MUX2X1 U12168 ( .B(n11230), .A(n11227), .S(n12585), .Y(n11241) );
  MUX2X1 U12169 ( .B(ram[874]), .A(ram[890]), .S(n12650), .Y(n11235) );
  MUX2X1 U12170 ( .B(ram[842]), .A(ram[858]), .S(n12669), .Y(n11234) );
  MUX2X1 U12171 ( .B(ram[810]), .A(ram[826]), .S(n12668), .Y(n11238) );
  MUX2X1 U12172 ( .B(ram[778]), .A(ram[794]), .S(n12663), .Y(n11237) );
  MUX2X1 U12173 ( .B(n11236), .A(n11233), .S(n12584), .Y(n11240) );
  MUX2X1 U12174 ( .B(ram[746]), .A(ram[762]), .S(n12636), .Y(n11244) );
  MUX2X1 U12175 ( .B(ram[714]), .A(ram[730]), .S(n12649), .Y(n11243) );
  MUX2X1 U12176 ( .B(ram[682]), .A(ram[698]), .S(n12637), .Y(n11247) );
  MUX2X1 U12177 ( .B(ram[650]), .A(ram[666]), .S(n12621), .Y(n11246) );
  MUX2X1 U12178 ( .B(n11245), .A(n11242), .S(n12583), .Y(n11256) );
  MUX2X1 U12179 ( .B(ram[618]), .A(ram[634]), .S(n12640), .Y(n11250) );
  MUX2X1 U12180 ( .B(ram[586]), .A(ram[602]), .S(mem_access_addr[0]), .Y(
        n11249) );
  MUX2X1 U12181 ( .B(ram[554]), .A(ram[570]), .S(n12639), .Y(n11253) );
  MUX2X1 U12182 ( .B(ram[522]), .A(ram[538]), .S(n12654), .Y(n11252) );
  MUX2X1 U12183 ( .B(n11251), .A(n11248), .S(n12576), .Y(n11255) );
  MUX2X1 U12184 ( .B(n11254), .A(n11239), .S(n12564), .Y(n11289) );
  MUX2X1 U12185 ( .B(ram[490]), .A(ram[506]), .S(n12648), .Y(n11259) );
  MUX2X1 U12186 ( .B(ram[458]), .A(ram[474]), .S(n12670), .Y(n11258) );
  MUX2X1 U12187 ( .B(ram[426]), .A(ram[442]), .S(n12648), .Y(n11262) );
  MUX2X1 U12188 ( .B(ram[394]), .A(ram[410]), .S(n12623), .Y(n11261) );
  MUX2X1 U12189 ( .B(n11260), .A(n11257), .S(n12579), .Y(n11271) );
  MUX2X1 U12190 ( .B(ram[362]), .A(ram[378]), .S(n12667), .Y(n11265) );
  MUX2X1 U12191 ( .B(ram[330]), .A(ram[346]), .S(n12623), .Y(n11264) );
  MUX2X1 U12192 ( .B(ram[298]), .A(ram[314]), .S(n12677), .Y(n11268) );
  MUX2X1 U12193 ( .B(ram[266]), .A(ram[282]), .S(n12622), .Y(n11267) );
  MUX2X1 U12194 ( .B(n11266), .A(n11263), .S(n12581), .Y(n11270) );
  MUX2X1 U12195 ( .B(ram[234]), .A(ram[250]), .S(n12661), .Y(n11274) );
  MUX2X1 U12196 ( .B(ram[202]), .A(ram[218]), .S(n12672), .Y(n11273) );
  MUX2X1 U12197 ( .B(ram[170]), .A(ram[186]), .S(n12639), .Y(n11277) );
  MUX2X1 U12198 ( .B(ram[138]), .A(ram[154]), .S(n12665), .Y(n11276) );
  MUX2X1 U12199 ( .B(n11275), .A(n11272), .S(n12582), .Y(n11286) );
  MUX2X1 U12200 ( .B(ram[106]), .A(ram[122]), .S(n12669), .Y(n11280) );
  MUX2X1 U12201 ( .B(ram[74]), .A(ram[90]), .S(n12661), .Y(n11279) );
  MUX2X1 U12202 ( .B(ram[42]), .A(ram[58]), .S(n12643), .Y(n11283) );
  MUX2X1 U12203 ( .B(ram[10]), .A(ram[26]), .S(n12644), .Y(n11282) );
  MUX2X1 U12204 ( .B(n11281), .A(n11278), .S(n12578), .Y(n11285) );
  MUX2X1 U12205 ( .B(n11284), .A(n11269), .S(n12565), .Y(n11288) );
  MUX2X1 U12206 ( .B(n11287), .A(n11224), .S(mem_access_addr[6]), .Y(n11290)
         );
  MUX2X1 U12207 ( .B(ram[4075]), .A(ram[4091]), .S(n12675), .Y(n11294) );
  MUX2X1 U12208 ( .B(ram[4043]), .A(ram[4059]), .S(n12636), .Y(n11293) );
  MUX2X1 U12209 ( .B(ram[4011]), .A(ram[4027]), .S(n12636), .Y(n11297) );
  MUX2X1 U12210 ( .B(ram[3979]), .A(ram[3995]), .S(n12647), .Y(n11296) );
  MUX2X1 U12211 ( .B(n11295), .A(n11292), .S(n12577), .Y(n11306) );
  MUX2X1 U12212 ( .B(ram[3947]), .A(ram[3963]), .S(n12660), .Y(n11300) );
  MUX2X1 U12213 ( .B(ram[3915]), .A(ram[3931]), .S(n12631), .Y(n11299) );
  MUX2X1 U12214 ( .B(ram[3883]), .A(ram[3899]), .S(n12677), .Y(n11303) );
  MUX2X1 U12215 ( .B(ram[3851]), .A(ram[3867]), .S(n12672), .Y(n11302) );
  MUX2X1 U12216 ( .B(n11301), .A(n11298), .S(n12577), .Y(n11305) );
  MUX2X1 U12217 ( .B(ram[3819]), .A(ram[3835]), .S(n12674), .Y(n11309) );
  MUX2X1 U12218 ( .B(ram[3787]), .A(ram[3803]), .S(n12667), .Y(n11308) );
  MUX2X1 U12219 ( .B(ram[3755]), .A(ram[3771]), .S(n12680), .Y(n11312) );
  MUX2X1 U12220 ( .B(ram[3723]), .A(ram[3739]), .S(n12666), .Y(n11311) );
  MUX2X1 U12221 ( .B(n11310), .A(n11307), .S(n12582), .Y(n11321) );
  MUX2X1 U12222 ( .B(ram[3691]), .A(ram[3707]), .S(n12627), .Y(n11315) );
  MUX2X1 U12223 ( .B(ram[3659]), .A(ram[3675]), .S(n12632), .Y(n11314) );
  MUX2X1 U12224 ( .B(ram[3627]), .A(ram[3643]), .S(n12627), .Y(n11318) );
  MUX2X1 U12225 ( .B(ram[3595]), .A(ram[3611]), .S(n12633), .Y(n11317) );
  MUX2X1 U12226 ( .B(n11316), .A(n11313), .S(n12580), .Y(n11320) );
  MUX2X1 U12227 ( .B(n11319), .A(n11304), .S(n12564), .Y(n11354) );
  MUX2X1 U12228 ( .B(ram[3563]), .A(ram[3579]), .S(n12649), .Y(n11324) );
  MUX2X1 U12229 ( .B(ram[3531]), .A(ram[3547]), .S(n12630), .Y(n11323) );
  MUX2X1 U12230 ( .B(ram[3499]), .A(ram[3515]), .S(n12639), .Y(n11327) );
  MUX2X1 U12231 ( .B(ram[3467]), .A(ram[3483]), .S(n12678), .Y(n11326) );
  MUX2X1 U12232 ( .B(n11325), .A(n11322), .S(n12581), .Y(n11336) );
  MUX2X1 U12233 ( .B(ram[3435]), .A(ram[3451]), .S(n12675), .Y(n11330) );
  MUX2X1 U12234 ( .B(ram[3403]), .A(ram[3419]), .S(n12680), .Y(n11329) );
  MUX2X1 U12235 ( .B(ram[3371]), .A(ram[3387]), .S(n12635), .Y(n11333) );
  MUX2X1 U12236 ( .B(ram[3339]), .A(ram[3355]), .S(n12673), .Y(n11332) );
  MUX2X1 U12237 ( .B(n11331), .A(n11328), .S(n12576), .Y(n11335) );
  MUX2X1 U12238 ( .B(ram[3307]), .A(ram[3323]), .S(n12642), .Y(n11339) );
  MUX2X1 U12239 ( .B(ram[3275]), .A(ram[3291]), .S(n12634), .Y(n11338) );
  MUX2X1 U12240 ( .B(ram[3243]), .A(ram[3259]), .S(n12654), .Y(n11342) );
  MUX2X1 U12241 ( .B(ram[3211]), .A(ram[3227]), .S(n12651), .Y(n11341) );
  MUX2X1 U12242 ( .B(n11340), .A(n11337), .S(n12583), .Y(n11351) );
  MUX2X1 U12243 ( .B(ram[3179]), .A(ram[3195]), .S(n12624), .Y(n11345) );
  MUX2X1 U12244 ( .B(ram[3147]), .A(ram[3163]), .S(n12641), .Y(n11344) );
  MUX2X1 U12245 ( .B(ram[3115]), .A(ram[3131]), .S(n12667), .Y(n11348) );
  MUX2X1 U12246 ( .B(ram[3083]), .A(ram[3099]), .S(n12649), .Y(n11347) );
  MUX2X1 U12247 ( .B(n11346), .A(n11343), .S(n12588), .Y(n11350) );
  MUX2X1 U12248 ( .B(n11349), .A(n11334), .S(n12564), .Y(n11353) );
  MUX2X1 U12249 ( .B(ram[3051]), .A(ram[3067]), .S(n12650), .Y(n11357) );
  MUX2X1 U12250 ( .B(ram[3019]), .A(ram[3035]), .S(n12653), .Y(n11356) );
  MUX2X1 U12251 ( .B(ram[2987]), .A(ram[3003]), .S(n12632), .Y(n11360) );
  MUX2X1 U12252 ( .B(ram[2955]), .A(ram[2971]), .S(n12671), .Y(n11359) );
  MUX2X1 U12253 ( .B(n11358), .A(n11355), .S(n12579), .Y(n11369) );
  MUX2X1 U12254 ( .B(ram[2923]), .A(ram[2939]), .S(n12652), .Y(n11363) );
  MUX2X1 U12255 ( .B(ram[2891]), .A(ram[2907]), .S(n12677), .Y(n11362) );
  MUX2X1 U12256 ( .B(ram[2859]), .A(ram[2875]), .S(n12642), .Y(n11366) );
  MUX2X1 U12257 ( .B(ram[2827]), .A(ram[2843]), .S(n12670), .Y(n11365) );
  MUX2X1 U12258 ( .B(n11364), .A(n11361), .S(n12584), .Y(n11368) );
  MUX2X1 U12259 ( .B(ram[2795]), .A(ram[2811]), .S(n12667), .Y(n11372) );
  MUX2X1 U12260 ( .B(ram[2763]), .A(ram[2779]), .S(n12629), .Y(n11371) );
  MUX2X1 U12261 ( .B(ram[2731]), .A(ram[2747]), .S(n12634), .Y(n11375) );
  MUX2X1 U12262 ( .B(ram[2699]), .A(ram[2715]), .S(n12628), .Y(n11374) );
  MUX2X1 U12263 ( .B(n11373), .A(n11370), .S(n12589), .Y(n11384) );
  MUX2X1 U12264 ( .B(ram[2667]), .A(ram[2683]), .S(n12649), .Y(n11378) );
  MUX2X1 U12265 ( .B(ram[2635]), .A(ram[2651]), .S(n12621), .Y(n11377) );
  MUX2X1 U12266 ( .B(ram[2603]), .A(ram[2619]), .S(n12638), .Y(n11381) );
  MUX2X1 U12267 ( .B(ram[2571]), .A(ram[2587]), .S(n12666), .Y(n11380) );
  MUX2X1 U12268 ( .B(n11379), .A(n11376), .S(n12585), .Y(n11383) );
  MUX2X1 U12269 ( .B(n11382), .A(n11367), .S(n12564), .Y(n11417) );
  MUX2X1 U12270 ( .B(ram[2539]), .A(ram[2555]), .S(n12642), .Y(n11387) );
  MUX2X1 U12271 ( .B(ram[2507]), .A(ram[2523]), .S(n12643), .Y(n11386) );
  MUX2X1 U12272 ( .B(ram[2475]), .A(ram[2491]), .S(n12664), .Y(n11390) );
  MUX2X1 U12273 ( .B(ram[2443]), .A(ram[2459]), .S(n12634), .Y(n11389) );
  MUX2X1 U12274 ( .B(n11388), .A(n11385), .S(n12578), .Y(n11399) );
  MUX2X1 U12275 ( .B(ram[2411]), .A(ram[2427]), .S(n12647), .Y(n11393) );
  MUX2X1 U12276 ( .B(ram[2379]), .A(ram[2395]), .S(n12638), .Y(n11392) );
  MUX2X1 U12277 ( .B(ram[2347]), .A(ram[2363]), .S(n12641), .Y(n11396) );
  MUX2X1 U12278 ( .B(ram[2315]), .A(ram[2331]), .S(n12671), .Y(n11395) );
  MUX2X1 U12279 ( .B(n11394), .A(n11391), .S(n12587), .Y(n11398) );
  MUX2X1 U12280 ( .B(ram[2283]), .A(ram[2299]), .S(n12625), .Y(n11402) );
  MUX2X1 U12281 ( .B(ram[2251]), .A(ram[2267]), .S(n12665), .Y(n11401) );
  MUX2X1 U12282 ( .B(ram[2219]), .A(ram[2235]), .S(n12632), .Y(n11405) );
  MUX2X1 U12283 ( .B(ram[2187]), .A(ram[2203]), .S(n12662), .Y(n11404) );
  MUX2X1 U12284 ( .B(n11403), .A(n11400), .S(n12582), .Y(n11414) );
  MUX2X1 U12285 ( .B(ram[2155]), .A(ram[2171]), .S(n12676), .Y(n11408) );
  MUX2X1 U12286 ( .B(ram[2123]), .A(ram[2139]), .S(n12645), .Y(n11407) );
  MUX2X1 U12287 ( .B(ram[2091]), .A(ram[2107]), .S(n12668), .Y(n11411) );
  MUX2X1 U12288 ( .B(ram[2059]), .A(ram[2075]), .S(n12658), .Y(n11410) );
  MUX2X1 U12289 ( .B(n11409), .A(n11406), .S(n12589), .Y(n11413) );
  MUX2X1 U12290 ( .B(n11412), .A(n11397), .S(n12564), .Y(n11416) );
  MUX2X1 U12291 ( .B(n11415), .A(n11352), .S(mem_access_addr[6]), .Y(n11545)
         );
  MUX2X1 U12292 ( .B(ram[2027]), .A(ram[2043]), .S(n12625), .Y(n11420) );
  MUX2X1 U12293 ( .B(ram[1995]), .A(ram[2011]), .S(n12635), .Y(n11419) );
  MUX2X1 U12294 ( .B(ram[1963]), .A(ram[1979]), .S(n12668), .Y(n11423) );
  MUX2X1 U12295 ( .B(ram[1931]), .A(ram[1947]), .S(n12682), .Y(n11422) );
  MUX2X1 U12296 ( .B(n11421), .A(n11418), .S(n12580), .Y(n11432) );
  MUX2X1 U12297 ( .B(ram[1899]), .A(ram[1915]), .S(n12638), .Y(n11426) );
  MUX2X1 U12298 ( .B(ram[1867]), .A(ram[1883]), .S(n12653), .Y(n11425) );
  MUX2X1 U12299 ( .B(ram[1835]), .A(ram[1851]), .S(n12674), .Y(n11429) );
  MUX2X1 U12300 ( .B(ram[1803]), .A(ram[1819]), .S(n12669), .Y(n11428) );
  MUX2X1 U12301 ( .B(n11427), .A(n11424), .S(n12584), .Y(n11431) );
  MUX2X1 U12302 ( .B(ram[1771]), .A(ram[1787]), .S(n12644), .Y(n11435) );
  MUX2X1 U12303 ( .B(ram[1739]), .A(ram[1755]), .S(n12661), .Y(n11434) );
  MUX2X1 U12304 ( .B(ram[1707]), .A(ram[1723]), .S(n12649), .Y(n11438) );
  MUX2X1 U12305 ( .B(ram[1675]), .A(ram[1691]), .S(n12623), .Y(n11437) );
  MUX2X1 U12306 ( .B(n11436), .A(n11433), .S(n12580), .Y(n11447) );
  MUX2X1 U12307 ( .B(ram[1643]), .A(ram[1659]), .S(n12627), .Y(n11441) );
  MUX2X1 U12308 ( .B(ram[1611]), .A(ram[1627]), .S(n12653), .Y(n11440) );
  MUX2X1 U12309 ( .B(ram[1579]), .A(ram[1595]), .S(n12651), .Y(n11444) );
  MUX2X1 U12310 ( .B(ram[1547]), .A(ram[1563]), .S(n12626), .Y(n11443) );
  MUX2X1 U12311 ( .B(n11442), .A(n11439), .S(n12581), .Y(n11446) );
  MUX2X1 U12312 ( .B(n11445), .A(n11430), .S(n12565), .Y(n11480) );
  MUX2X1 U12313 ( .B(ram[1515]), .A(ram[1531]), .S(n12659), .Y(n11450) );
  MUX2X1 U12314 ( .B(ram[1483]), .A(ram[1499]), .S(n12662), .Y(n11449) );
  MUX2X1 U12315 ( .B(ram[1451]), .A(ram[1467]), .S(n12633), .Y(n11453) );
  MUX2X1 U12316 ( .B(ram[1419]), .A(ram[1435]), .S(n12652), .Y(n11452) );
  MUX2X1 U12317 ( .B(n11451), .A(n11448), .S(n12577), .Y(n11462) );
  MUX2X1 U12318 ( .B(ram[1387]), .A(ram[1403]), .S(n12622), .Y(n11456) );
  MUX2X1 U12319 ( .B(ram[1355]), .A(ram[1371]), .S(n12642), .Y(n11455) );
  MUX2X1 U12320 ( .B(ram[1323]), .A(ram[1339]), .S(n12634), .Y(n11459) );
  MUX2X1 U12321 ( .B(ram[1291]), .A(ram[1307]), .S(n12624), .Y(n11458) );
  MUX2X1 U12322 ( .B(n11457), .A(n11454), .S(n12583), .Y(n11461) );
  MUX2X1 U12323 ( .B(ram[1259]), .A(ram[1275]), .S(n12631), .Y(n11465) );
  MUX2X1 U12324 ( .B(ram[1227]), .A(ram[1243]), .S(n12623), .Y(n11464) );
  MUX2X1 U12325 ( .B(ram[1195]), .A(ram[1211]), .S(n12624), .Y(n11468) );
  MUX2X1 U12326 ( .B(ram[1163]), .A(ram[1179]), .S(n12637), .Y(n11467) );
  MUX2X1 U12327 ( .B(n11466), .A(n11463), .S(n12582), .Y(n11477) );
  MUX2X1 U12328 ( .B(ram[1131]), .A(ram[1147]), .S(n12664), .Y(n11471) );
  MUX2X1 U12329 ( .B(ram[1099]), .A(ram[1115]), .S(n12683), .Y(n11470) );
  MUX2X1 U12330 ( .B(ram[1067]), .A(ram[1083]), .S(n12633), .Y(n11474) );
  MUX2X1 U12331 ( .B(ram[1035]), .A(ram[1051]), .S(n12622), .Y(n11473) );
  MUX2X1 U12332 ( .B(n11472), .A(n11469), .S(n12581), .Y(n11476) );
  MUX2X1 U12333 ( .B(n11475), .A(n11460), .S(n12565), .Y(n11479) );
  MUX2X1 U12334 ( .B(ram[1003]), .A(ram[1019]), .S(n12634), .Y(n11483) );
  MUX2X1 U12335 ( .B(ram[971]), .A(ram[987]), .S(n12644), .Y(n11482) );
  MUX2X1 U12336 ( .B(ram[939]), .A(ram[955]), .S(n12629), .Y(n11486) );
  MUX2X1 U12337 ( .B(ram[907]), .A(ram[923]), .S(n12660), .Y(n11485) );
  MUX2X1 U12338 ( .B(n11484), .A(n11481), .S(n12585), .Y(n11495) );
  MUX2X1 U12339 ( .B(ram[875]), .A(ram[891]), .S(n12672), .Y(n11489) );
  MUX2X1 U12340 ( .B(ram[843]), .A(ram[859]), .S(n12668), .Y(n11488) );
  MUX2X1 U12341 ( .B(ram[811]), .A(ram[827]), .S(n12674), .Y(n11492) );
  MUX2X1 U12342 ( .B(ram[779]), .A(ram[795]), .S(n12655), .Y(n11491) );
  MUX2X1 U12343 ( .B(n11490), .A(n11487), .S(n12579), .Y(n11494) );
  MUX2X1 U12344 ( .B(ram[747]), .A(ram[763]), .S(n12621), .Y(n11498) );
  MUX2X1 U12345 ( .B(ram[715]), .A(ram[731]), .S(n12659), .Y(n11497) );
  MUX2X1 U12346 ( .B(ram[683]), .A(ram[699]), .S(n12636), .Y(n11501) );
  MUX2X1 U12347 ( .B(ram[651]), .A(ram[667]), .S(n12650), .Y(n11500) );
  MUX2X1 U12348 ( .B(n11499), .A(n11496), .S(n12582), .Y(n11510) );
  MUX2X1 U12349 ( .B(ram[619]), .A(ram[635]), .S(n12636), .Y(n11504) );
  MUX2X1 U12350 ( .B(ram[587]), .A(ram[603]), .S(n12641), .Y(n11503) );
  MUX2X1 U12351 ( .B(ram[555]), .A(ram[571]), .S(n12670), .Y(n11507) );
  MUX2X1 U12352 ( .B(ram[523]), .A(ram[539]), .S(n12632), .Y(n11506) );
  MUX2X1 U12353 ( .B(n11505), .A(n11502), .S(n12578), .Y(n11509) );
  MUX2X1 U12354 ( .B(n11508), .A(n11493), .S(n12565), .Y(n11543) );
  MUX2X1 U12355 ( .B(ram[491]), .A(ram[507]), .S(n12641), .Y(n11513) );
  MUX2X1 U12356 ( .B(ram[459]), .A(ram[475]), .S(n12647), .Y(n11512) );
  MUX2X1 U12357 ( .B(ram[427]), .A(ram[443]), .S(n12621), .Y(n11516) );
  MUX2X1 U12358 ( .B(ram[395]), .A(ram[411]), .S(n12637), .Y(n11515) );
  MUX2X1 U12359 ( .B(n11514), .A(n11511), .S(n12585), .Y(n11525) );
  MUX2X1 U12360 ( .B(ram[363]), .A(ram[379]), .S(n12626), .Y(n11519) );
  MUX2X1 U12361 ( .B(ram[331]), .A(ram[347]), .S(n12652), .Y(n11518) );
  MUX2X1 U12362 ( .B(ram[299]), .A(ram[315]), .S(n12663), .Y(n11522) );
  MUX2X1 U12363 ( .B(ram[267]), .A(ram[283]), .S(n12625), .Y(n11521) );
  MUX2X1 U12364 ( .B(n11520), .A(n11517), .S(n12584), .Y(n11524) );
  MUX2X1 U12365 ( .B(ram[235]), .A(ram[251]), .S(n12662), .Y(n11528) );
  MUX2X1 U12366 ( .B(ram[203]), .A(ram[219]), .S(n12660), .Y(n11527) );
  MUX2X1 U12367 ( .B(ram[171]), .A(ram[187]), .S(n12681), .Y(n11531) );
  MUX2X1 U12368 ( .B(ram[139]), .A(ram[155]), .S(n12672), .Y(n11530) );
  MUX2X1 U12369 ( .B(n11529), .A(n11526), .S(n12576), .Y(n11540) );
  MUX2X1 U12370 ( .B(ram[107]), .A(ram[123]), .S(n12634), .Y(n11534) );
  MUX2X1 U12371 ( .B(ram[75]), .A(ram[91]), .S(n12646), .Y(n11533) );
  MUX2X1 U12372 ( .B(ram[43]), .A(ram[59]), .S(n12644), .Y(n11537) );
  MUX2X1 U12373 ( .B(ram[11]), .A(ram[27]), .S(n12630), .Y(n11536) );
  MUX2X1 U12374 ( .B(n11535), .A(n11532), .S(n12579), .Y(n11539) );
  MUX2X1 U12375 ( .B(n11538), .A(n11523), .S(n12565), .Y(n11542) );
  MUX2X1 U12376 ( .B(n11541), .A(n11478), .S(mem_access_addr[6]), .Y(n11544)
         );
  MUX2X1 U12377 ( .B(ram[4076]), .A(ram[4092]), .S(n12637), .Y(n11548) );
  MUX2X1 U12378 ( .B(ram[4044]), .A(ram[4060]), .S(n12658), .Y(n11547) );
  MUX2X1 U12379 ( .B(ram[4012]), .A(ram[4028]), .S(n12679), .Y(n11551) );
  MUX2X1 U12380 ( .B(ram[3980]), .A(ram[3996]), .S(n12661), .Y(n11550) );
  MUX2X1 U12381 ( .B(n11549), .A(n11546), .S(n12580), .Y(n11560) );
  MUX2X1 U12382 ( .B(ram[3948]), .A(ram[3964]), .S(n12676), .Y(n11554) );
  MUX2X1 U12383 ( .B(ram[3916]), .A(ram[3932]), .S(n12639), .Y(n11553) );
  MUX2X1 U12384 ( .B(ram[3884]), .A(ram[3900]), .S(n12651), .Y(n11557) );
  MUX2X1 U12385 ( .B(ram[3852]), .A(ram[3868]), .S(n12673), .Y(n11556) );
  MUX2X1 U12386 ( .B(n11555), .A(n11552), .S(n12577), .Y(n11559) );
  MUX2X1 U12387 ( .B(ram[3820]), .A(ram[3836]), .S(n12657), .Y(n11563) );
  MUX2X1 U12388 ( .B(ram[3788]), .A(ram[3804]), .S(n12664), .Y(n11562) );
  MUX2X1 U12389 ( .B(ram[3756]), .A(ram[3772]), .S(n12631), .Y(n11566) );
  MUX2X1 U12390 ( .B(ram[3724]), .A(ram[3740]), .S(n12656), .Y(n11565) );
  MUX2X1 U12391 ( .B(n11564), .A(n11561), .S(n12578), .Y(n11575) );
  MUX2X1 U12392 ( .B(ram[3692]), .A(ram[3708]), .S(n12677), .Y(n11569) );
  MUX2X1 U12393 ( .B(ram[3660]), .A(ram[3676]), .S(n12631), .Y(n11568) );
  MUX2X1 U12394 ( .B(ram[3628]), .A(ram[3644]), .S(n12646), .Y(n11572) );
  MUX2X1 U12395 ( .B(ram[3596]), .A(ram[3612]), .S(n12665), .Y(n11571) );
  MUX2X1 U12396 ( .B(n11570), .A(n11567), .S(n12584), .Y(n11574) );
  MUX2X1 U12397 ( .B(n11573), .A(n11558), .S(n12565), .Y(n11608) );
  MUX2X1 U12398 ( .B(ram[3564]), .A(ram[3580]), .S(n12628), .Y(n11578) );
  MUX2X1 U12399 ( .B(ram[3532]), .A(ram[3548]), .S(n12640), .Y(n11577) );
  MUX2X1 U12400 ( .B(ram[3500]), .A(ram[3516]), .S(n12678), .Y(n11581) );
  MUX2X1 U12401 ( .B(ram[3468]), .A(ram[3484]), .S(n12647), .Y(n11580) );
  MUX2X1 U12402 ( .B(n11579), .A(n11576), .S(n12580), .Y(n11590) );
  MUX2X1 U12403 ( .B(ram[3436]), .A(ram[3452]), .S(n12659), .Y(n11584) );
  MUX2X1 U12404 ( .B(ram[3404]), .A(ram[3420]), .S(n12680), .Y(n11583) );
  MUX2X1 U12405 ( .B(ram[3372]), .A(ram[3388]), .S(n12646), .Y(n11587) );
  MUX2X1 U12406 ( .B(ram[3340]), .A(ram[3356]), .S(n12677), .Y(n11586) );
  MUX2X1 U12407 ( .B(n11585), .A(n11582), .S(n12585), .Y(n11589) );
  MUX2X1 U12408 ( .B(ram[3308]), .A(ram[3324]), .S(n12664), .Y(n11593) );
  MUX2X1 U12409 ( .B(ram[3276]), .A(ram[3292]), .S(n12638), .Y(n11592) );
  MUX2X1 U12410 ( .B(ram[3244]), .A(ram[3260]), .S(n12639), .Y(n11596) );
  MUX2X1 U12411 ( .B(ram[3212]), .A(ram[3228]), .S(n12678), .Y(n11595) );
  MUX2X1 U12412 ( .B(n11594), .A(n11591), .S(n12581), .Y(n11605) );
  MUX2X1 U12413 ( .B(ram[3180]), .A(ram[3196]), .S(n12670), .Y(n11599) );
  MUX2X1 U12414 ( .B(ram[3148]), .A(ram[3164]), .S(n12678), .Y(n11598) );
  MUX2X1 U12415 ( .B(ram[3116]), .A(ram[3132]), .S(n12677), .Y(n11602) );
  MUX2X1 U12416 ( .B(ram[3084]), .A(ram[3100]), .S(n12666), .Y(n11601) );
  MUX2X1 U12417 ( .B(n11600), .A(n11597), .S(n12583), .Y(n11604) );
  MUX2X1 U12418 ( .B(n11603), .A(n11588), .S(n12565), .Y(n11607) );
  MUX2X1 U12419 ( .B(ram[3052]), .A(ram[3068]), .S(n12645), .Y(n11611) );
  MUX2X1 U12420 ( .B(ram[3020]), .A(ram[3036]), .S(n12625), .Y(n11610) );
  MUX2X1 U12421 ( .B(ram[2988]), .A(ram[3004]), .S(n12630), .Y(n11614) );
  MUX2X1 U12422 ( .B(ram[2956]), .A(ram[2972]), .S(n12671), .Y(n11613) );
  MUX2X1 U12423 ( .B(n11612), .A(n11609), .S(n12576), .Y(n11623) );
  MUX2X1 U12424 ( .B(ram[2924]), .A(ram[2940]), .S(n12638), .Y(n11617) );
  MUX2X1 U12425 ( .B(ram[2892]), .A(ram[2908]), .S(n12662), .Y(n11616) );
  MUX2X1 U12426 ( .B(ram[2860]), .A(ram[2876]), .S(n12636), .Y(n11620) );
  MUX2X1 U12427 ( .B(ram[2828]), .A(ram[2844]), .S(n12659), .Y(n11619) );
  MUX2X1 U12428 ( .B(n11618), .A(n11615), .S(n12576), .Y(n11622) );
  MUX2X1 U12429 ( .B(ram[2796]), .A(ram[2812]), .S(n12635), .Y(n11626) );
  MUX2X1 U12430 ( .B(ram[2764]), .A(ram[2780]), .S(n12652), .Y(n11625) );
  MUX2X1 U12431 ( .B(ram[2732]), .A(ram[2748]), .S(n12647), .Y(n11629) );
  MUX2X1 U12432 ( .B(ram[2700]), .A(ram[2716]), .S(n12634), .Y(n11628) );
  MUX2X1 U12433 ( .B(n11627), .A(n11624), .S(n12576), .Y(n11638) );
  MUX2X1 U12434 ( .B(ram[2668]), .A(ram[2684]), .S(n12645), .Y(n11632) );
  MUX2X1 U12435 ( .B(ram[2636]), .A(ram[2652]), .S(n12627), .Y(n11631) );
  MUX2X1 U12436 ( .B(ram[2604]), .A(ram[2620]), .S(n12647), .Y(n11635) );
  MUX2X1 U12437 ( .B(ram[2572]), .A(ram[2588]), .S(n12631), .Y(n11634) );
  MUX2X1 U12438 ( .B(n11633), .A(n11630), .S(n12576), .Y(n11637) );
  MUX2X1 U12439 ( .B(n11636), .A(n11621), .S(n12565), .Y(n11671) );
  MUX2X1 U12440 ( .B(ram[2540]), .A(ram[2556]), .S(n12673), .Y(n11641) );
  MUX2X1 U12441 ( .B(ram[2508]), .A(ram[2524]), .S(n12670), .Y(n11640) );
  MUX2X1 U12442 ( .B(ram[2476]), .A(ram[2492]), .S(n12646), .Y(n11644) );
  MUX2X1 U12443 ( .B(ram[2444]), .A(ram[2460]), .S(n12624), .Y(n11643) );
  MUX2X1 U12444 ( .B(n11642), .A(n11639), .S(n12576), .Y(n11653) );
  MUX2X1 U12445 ( .B(ram[2412]), .A(ram[2428]), .S(n12629), .Y(n11647) );
  MUX2X1 U12446 ( .B(ram[2380]), .A(ram[2396]), .S(n12637), .Y(n11646) );
  MUX2X1 U12447 ( .B(ram[2348]), .A(ram[2364]), .S(n12645), .Y(n11650) );
  MUX2X1 U12448 ( .B(ram[2316]), .A(ram[2332]), .S(n12666), .Y(n11649) );
  MUX2X1 U12449 ( .B(n11648), .A(n11645), .S(n12576), .Y(n11652) );
  MUX2X1 U12450 ( .B(ram[2284]), .A(ram[2300]), .S(n12637), .Y(n11656) );
  MUX2X1 U12451 ( .B(ram[2252]), .A(ram[2268]), .S(n12638), .Y(n11655) );
  MUX2X1 U12452 ( .B(ram[2220]), .A(ram[2236]), .S(n12638), .Y(n11659) );
  MUX2X1 U12453 ( .B(ram[2188]), .A(ram[2204]), .S(n12622), .Y(n11658) );
  MUX2X1 U12454 ( .B(n11657), .A(n11654), .S(n12576), .Y(n11668) );
  MUX2X1 U12455 ( .B(ram[2156]), .A(ram[2172]), .S(n12625), .Y(n11662) );
  MUX2X1 U12456 ( .B(ram[2124]), .A(ram[2140]), .S(n12624), .Y(n11661) );
  MUX2X1 U12457 ( .B(ram[2092]), .A(ram[2108]), .S(n12630), .Y(n11665) );
  MUX2X1 U12458 ( .B(ram[2060]), .A(ram[2076]), .S(n12623), .Y(n11664) );
  MUX2X1 U12459 ( .B(n11663), .A(n11660), .S(n12576), .Y(n11667) );
  MUX2X1 U12460 ( .B(n11666), .A(n11651), .S(n12565), .Y(n11670) );
  MUX2X1 U12461 ( .B(n11669), .A(n11606), .S(mem_access_addr[6]), .Y(n11799)
         );
  MUX2X1 U12462 ( .B(ram[2028]), .A(ram[2044]), .S(n12637), .Y(n11674) );
  MUX2X1 U12463 ( .B(ram[1996]), .A(ram[2012]), .S(n12641), .Y(n11673) );
  MUX2X1 U12464 ( .B(ram[1964]), .A(ram[1980]), .S(n12628), .Y(n11677) );
  MUX2X1 U12465 ( .B(ram[1932]), .A(ram[1948]), .S(n12656), .Y(n11676) );
  MUX2X1 U12466 ( .B(n11675), .A(n11672), .S(n12576), .Y(n11686) );
  MUX2X1 U12467 ( .B(ram[1900]), .A(ram[1916]), .S(n12623), .Y(n11680) );
  MUX2X1 U12468 ( .B(ram[1868]), .A(ram[1884]), .S(n12623), .Y(n11679) );
  MUX2X1 U12469 ( .B(ram[1836]), .A(ram[1852]), .S(n12623), .Y(n11683) );
  MUX2X1 U12470 ( .B(ram[1804]), .A(ram[1820]), .S(n12655), .Y(n11682) );
  MUX2X1 U12471 ( .B(n11681), .A(n11678), .S(n12576), .Y(n11685) );
  MUX2X1 U12472 ( .B(ram[1772]), .A(ram[1788]), .S(n12629), .Y(n11689) );
  MUX2X1 U12473 ( .B(ram[1740]), .A(ram[1756]), .S(n12624), .Y(n11688) );
  MUX2X1 U12474 ( .B(ram[1708]), .A(ram[1724]), .S(n12631), .Y(n11692) );
  MUX2X1 U12475 ( .B(ram[1676]), .A(ram[1692]), .S(n12631), .Y(n11691) );
  MUX2X1 U12476 ( .B(n11690), .A(n11687), .S(n12576), .Y(n11701) );
  MUX2X1 U12477 ( .B(ram[1644]), .A(ram[1660]), .S(n12622), .Y(n11695) );
  MUX2X1 U12478 ( .B(ram[1612]), .A(ram[1628]), .S(n12622), .Y(n11694) );
  MUX2X1 U12479 ( .B(ram[1580]), .A(ram[1596]), .S(n12622), .Y(n11698) );
  MUX2X1 U12480 ( .B(ram[1548]), .A(ram[1564]), .S(n12624), .Y(n11697) );
  MUX2X1 U12481 ( .B(n11696), .A(n11693), .S(n12576), .Y(n11700) );
  MUX2X1 U12482 ( .B(n11699), .A(n11684), .S(n12565), .Y(n11734) );
  MUX2X1 U12483 ( .B(ram[1516]), .A(ram[1532]), .S(n12683), .Y(n11704) );
  MUX2X1 U12484 ( .B(ram[1484]), .A(ram[1500]), .S(n12682), .Y(n11703) );
  MUX2X1 U12485 ( .B(ram[1452]), .A(ram[1468]), .S(n12670), .Y(n11707) );
  MUX2X1 U12486 ( .B(ram[1420]), .A(ram[1436]), .S(n12683), .Y(n11706) );
  MUX2X1 U12487 ( .B(n11705), .A(n11702), .S(n12577), .Y(n11716) );
  MUX2X1 U12488 ( .B(ram[1388]), .A(ram[1404]), .S(n12682), .Y(n11710) );
  MUX2X1 U12489 ( .B(ram[1356]), .A(ram[1372]), .S(n12682), .Y(n11709) );
  MUX2X1 U12490 ( .B(ram[1324]), .A(ram[1340]), .S(n12621), .Y(n11713) );
  MUX2X1 U12491 ( .B(ram[1292]), .A(ram[1308]), .S(n12683), .Y(n11712) );
  MUX2X1 U12492 ( .B(n11711), .A(n11708), .S(n12577), .Y(n11715) );
  MUX2X1 U12493 ( .B(ram[1260]), .A(ram[1276]), .S(n12628), .Y(n11719) );
  MUX2X1 U12494 ( .B(ram[1228]), .A(ram[1244]), .S(n12643), .Y(n11718) );
  MUX2X1 U12495 ( .B(ram[1196]), .A(ram[1212]), .S(n12622), .Y(n11722) );
  MUX2X1 U12496 ( .B(ram[1164]), .A(ram[1180]), .S(n12667), .Y(n11721) );
  MUX2X1 U12497 ( .B(n11720), .A(n11717), .S(n12577), .Y(n11731) );
  MUX2X1 U12498 ( .B(ram[1132]), .A(ram[1148]), .S(n12648), .Y(n11725) );
  MUX2X1 U12499 ( .B(ram[1100]), .A(ram[1116]), .S(n12648), .Y(n11724) );
  MUX2X1 U12500 ( .B(ram[1068]), .A(ram[1084]), .S(n12648), .Y(n11728) );
  MUX2X1 U12501 ( .B(ram[1036]), .A(ram[1052]), .S(n12648), .Y(n11727) );
  MUX2X1 U12502 ( .B(n11726), .A(n11723), .S(n12577), .Y(n11730) );
  MUX2X1 U12503 ( .B(n11729), .A(n11714), .S(n12565), .Y(n11733) );
  MUX2X1 U12504 ( .B(ram[1004]), .A(ram[1020]), .S(n12648), .Y(n11737) );
  MUX2X1 U12505 ( .B(ram[972]), .A(ram[988]), .S(n12648), .Y(n11736) );
  MUX2X1 U12506 ( .B(ram[940]), .A(ram[956]), .S(n12648), .Y(n11740) );
  MUX2X1 U12507 ( .B(ram[908]), .A(ram[924]), .S(n12648), .Y(n11739) );
  MUX2X1 U12508 ( .B(n11738), .A(n11735), .S(n12577), .Y(n11749) );
  MUX2X1 U12509 ( .B(ram[876]), .A(ram[892]), .S(n12648), .Y(n11743) );
  MUX2X1 U12510 ( .B(ram[844]), .A(ram[860]), .S(n12648), .Y(n11742) );
  MUX2X1 U12511 ( .B(ram[812]), .A(ram[828]), .S(n12648), .Y(n11746) );
  MUX2X1 U12512 ( .B(ram[780]), .A(ram[796]), .S(n12648), .Y(n11745) );
  MUX2X1 U12513 ( .B(n11744), .A(n11741), .S(n12577), .Y(n11748) );
  MUX2X1 U12514 ( .B(ram[748]), .A(ram[764]), .S(n12622), .Y(n11752) );
  MUX2X1 U12515 ( .B(ram[716]), .A(ram[732]), .S(n12629), .Y(n11751) );
  MUX2X1 U12516 ( .B(ram[684]), .A(ram[700]), .S(n12661), .Y(n11755) );
  MUX2X1 U12517 ( .B(ram[652]), .A(ram[668]), .S(n12625), .Y(n11754) );
  MUX2X1 U12518 ( .B(n11753), .A(n11750), .S(n12577), .Y(n11764) );
  MUX2X1 U12519 ( .B(ram[620]), .A(ram[636]), .S(n12672), .Y(n11758) );
  MUX2X1 U12520 ( .B(ram[588]), .A(ram[604]), .S(n12683), .Y(n11757) );
  MUX2X1 U12521 ( .B(ram[556]), .A(ram[572]), .S(n12669), .Y(n11761) );
  MUX2X1 U12522 ( .B(ram[524]), .A(ram[540]), .S(n12639), .Y(n11760) );
  MUX2X1 U12523 ( .B(n11759), .A(n11756), .S(n12577), .Y(n11763) );
  MUX2X1 U12524 ( .B(n11762), .A(n11747), .S(n12565), .Y(n11797) );
  MUX2X1 U12525 ( .B(ram[492]), .A(ram[508]), .S(n12683), .Y(n11767) );
  MUX2X1 U12526 ( .B(ram[460]), .A(ram[476]), .S(n12682), .Y(n11766) );
  MUX2X1 U12527 ( .B(ram[428]), .A(ram[444]), .S(n12671), .Y(n11770) );
  MUX2X1 U12528 ( .B(ram[396]), .A(ram[412]), .S(n12682), .Y(n11769) );
  MUX2X1 U12529 ( .B(n11768), .A(n11765), .S(n12577), .Y(n11779) );
  MUX2X1 U12530 ( .B(ram[364]), .A(ram[380]), .S(n12649), .Y(n11773) );
  MUX2X1 U12531 ( .B(ram[332]), .A(ram[348]), .S(n12649), .Y(n11772) );
  MUX2X1 U12532 ( .B(ram[300]), .A(ram[316]), .S(n12649), .Y(n11776) );
  MUX2X1 U12533 ( .B(ram[268]), .A(ram[284]), .S(n12649), .Y(n11775) );
  MUX2X1 U12534 ( .B(n11774), .A(n11771), .S(n12577), .Y(n11778) );
  MUX2X1 U12535 ( .B(ram[236]), .A(ram[252]), .S(n12649), .Y(n11782) );
  MUX2X1 U12536 ( .B(ram[204]), .A(ram[220]), .S(n12649), .Y(n11781) );
  MUX2X1 U12537 ( .B(ram[172]), .A(ram[188]), .S(n12649), .Y(n11785) );
  MUX2X1 U12538 ( .B(ram[140]), .A(ram[156]), .S(n12649), .Y(n11784) );
  MUX2X1 U12539 ( .B(n11783), .A(n11780), .S(n12577), .Y(n11794) );
  MUX2X1 U12540 ( .B(ram[108]), .A(ram[124]), .S(n12649), .Y(n11788) );
  MUX2X1 U12541 ( .B(ram[76]), .A(ram[92]), .S(n12649), .Y(n11787) );
  MUX2X1 U12542 ( .B(ram[44]), .A(ram[60]), .S(n12649), .Y(n11791) );
  MUX2X1 U12543 ( .B(ram[12]), .A(ram[28]), .S(n12649), .Y(n11790) );
  MUX2X1 U12544 ( .B(n11789), .A(n11786), .S(n12577), .Y(n11793) );
  MUX2X1 U12545 ( .B(n11792), .A(n11777), .S(n12565), .Y(n11796) );
  MUX2X1 U12546 ( .B(n11795), .A(n11732), .S(mem_access_addr[6]), .Y(n11798)
         );
  MUX2X1 U12547 ( .B(ram[4077]), .A(ram[4093]), .S(n12650), .Y(n11802) );
  MUX2X1 U12548 ( .B(ram[4045]), .A(ram[4061]), .S(n12650), .Y(n11801) );
  MUX2X1 U12549 ( .B(ram[4013]), .A(ram[4029]), .S(n12650), .Y(n11805) );
  MUX2X1 U12550 ( .B(ram[3981]), .A(ram[3997]), .S(n12650), .Y(n11804) );
  MUX2X1 U12551 ( .B(n11803), .A(n11800), .S(n12578), .Y(n11814) );
  MUX2X1 U12552 ( .B(ram[3949]), .A(ram[3965]), .S(n12650), .Y(n11808) );
  MUX2X1 U12553 ( .B(ram[3917]), .A(ram[3933]), .S(n12650), .Y(n11807) );
  MUX2X1 U12554 ( .B(ram[3885]), .A(ram[3901]), .S(n12650), .Y(n11811) );
  MUX2X1 U12555 ( .B(ram[3853]), .A(ram[3869]), .S(n12650), .Y(n11810) );
  MUX2X1 U12556 ( .B(n11809), .A(n11806), .S(n12578), .Y(n11813) );
  MUX2X1 U12557 ( .B(ram[3821]), .A(ram[3837]), .S(n12650), .Y(n11817) );
  MUX2X1 U12558 ( .B(ram[3789]), .A(ram[3805]), .S(n12650), .Y(n11816) );
  MUX2X1 U12559 ( .B(ram[3757]), .A(ram[3773]), .S(n12650), .Y(n11820) );
  MUX2X1 U12560 ( .B(ram[3725]), .A(ram[3741]), .S(n12650), .Y(n11819) );
  MUX2X1 U12561 ( .B(n11818), .A(n11815), .S(n12578), .Y(n11829) );
  MUX2X1 U12562 ( .B(ram[3693]), .A(ram[3709]), .S(n12651), .Y(n11823) );
  MUX2X1 U12563 ( .B(ram[3661]), .A(ram[3677]), .S(n12651), .Y(n11822) );
  MUX2X1 U12564 ( .B(ram[3629]), .A(ram[3645]), .S(n12651), .Y(n11826) );
  MUX2X1 U12565 ( .B(ram[3597]), .A(ram[3613]), .S(n12651), .Y(n11825) );
  MUX2X1 U12566 ( .B(n11824), .A(n11821), .S(n12578), .Y(n11828) );
  MUX2X1 U12567 ( .B(n11827), .A(n11812), .S(n12566), .Y(n11862) );
  MUX2X1 U12568 ( .B(ram[3565]), .A(ram[3581]), .S(n12651), .Y(n11832) );
  MUX2X1 U12569 ( .B(ram[3533]), .A(ram[3549]), .S(n12651), .Y(n11831) );
  MUX2X1 U12570 ( .B(ram[3501]), .A(ram[3517]), .S(n12651), .Y(n11835) );
  MUX2X1 U12571 ( .B(ram[3469]), .A(ram[3485]), .S(n12651), .Y(n11834) );
  MUX2X1 U12572 ( .B(n11833), .A(n11830), .S(n12578), .Y(n11844) );
  MUX2X1 U12573 ( .B(ram[3437]), .A(ram[3453]), .S(n12651), .Y(n11838) );
  MUX2X1 U12574 ( .B(ram[3405]), .A(ram[3421]), .S(n12651), .Y(n11837) );
  MUX2X1 U12575 ( .B(ram[3373]), .A(ram[3389]), .S(n12651), .Y(n11841) );
  MUX2X1 U12576 ( .B(ram[3341]), .A(ram[3357]), .S(n12651), .Y(n11840) );
  MUX2X1 U12577 ( .B(n11839), .A(n11836), .S(n12578), .Y(n11843) );
  MUX2X1 U12578 ( .B(ram[3309]), .A(ram[3325]), .S(n12652), .Y(n11847) );
  MUX2X1 U12579 ( .B(ram[3277]), .A(ram[3293]), .S(n12652), .Y(n11846) );
  MUX2X1 U12580 ( .B(ram[3245]), .A(ram[3261]), .S(n12652), .Y(n11850) );
  MUX2X1 U12581 ( .B(ram[3213]), .A(ram[3229]), .S(n12652), .Y(n11849) );
  MUX2X1 U12582 ( .B(n11848), .A(n11845), .S(n12578), .Y(n11859) );
  MUX2X1 U12583 ( .B(ram[3181]), .A(ram[3197]), .S(n12652), .Y(n11853) );
  MUX2X1 U12584 ( .B(ram[3149]), .A(ram[3165]), .S(n12652), .Y(n11852) );
  MUX2X1 U12585 ( .B(ram[3117]), .A(ram[3133]), .S(n12652), .Y(n11856) );
  MUX2X1 U12586 ( .B(ram[3085]), .A(ram[3101]), .S(n12652), .Y(n11855) );
  MUX2X1 U12587 ( .B(n11854), .A(n11851), .S(n12578), .Y(n11858) );
  MUX2X1 U12588 ( .B(n11857), .A(n11842), .S(n12566), .Y(n11861) );
  MUX2X1 U12589 ( .B(ram[3053]), .A(ram[3069]), .S(n12652), .Y(n11865) );
  MUX2X1 U12590 ( .B(ram[3021]), .A(ram[3037]), .S(n12652), .Y(n11864) );
  MUX2X1 U12591 ( .B(ram[2989]), .A(ram[3005]), .S(n12652), .Y(n11868) );
  MUX2X1 U12592 ( .B(ram[2957]), .A(ram[2973]), .S(n12652), .Y(n11867) );
  MUX2X1 U12593 ( .B(n11866), .A(n11863), .S(n12578), .Y(n11877) );
  MUX2X1 U12594 ( .B(ram[2925]), .A(ram[2941]), .S(n12653), .Y(n11871) );
  MUX2X1 U12595 ( .B(ram[2893]), .A(ram[2909]), .S(n12653), .Y(n11870) );
  MUX2X1 U12596 ( .B(ram[2861]), .A(ram[2877]), .S(n12653), .Y(n11874) );
  MUX2X1 U12597 ( .B(ram[2829]), .A(ram[2845]), .S(n12653), .Y(n11873) );
  MUX2X1 U12598 ( .B(n11872), .A(n11869), .S(n12578), .Y(n11876) );
  MUX2X1 U12599 ( .B(ram[2797]), .A(ram[2813]), .S(n12653), .Y(n11880) );
  MUX2X1 U12600 ( .B(ram[2765]), .A(ram[2781]), .S(n12653), .Y(n11879) );
  MUX2X1 U12601 ( .B(ram[2733]), .A(ram[2749]), .S(n12653), .Y(n11883) );
  MUX2X1 U12602 ( .B(ram[2701]), .A(ram[2717]), .S(n12653), .Y(n11882) );
  MUX2X1 U12603 ( .B(n11881), .A(n11878), .S(n12578), .Y(n11892) );
  MUX2X1 U12604 ( .B(ram[2669]), .A(ram[2685]), .S(n12653), .Y(n11886) );
  MUX2X1 U12605 ( .B(ram[2637]), .A(ram[2653]), .S(n12653), .Y(n11885) );
  MUX2X1 U12606 ( .B(ram[2605]), .A(ram[2621]), .S(n12653), .Y(n11889) );
  MUX2X1 U12607 ( .B(ram[2573]), .A(ram[2589]), .S(n12653), .Y(n11888) );
  MUX2X1 U12608 ( .B(n11887), .A(n11884), .S(n12578), .Y(n11891) );
  MUX2X1 U12609 ( .B(n11890), .A(n11875), .S(n12566), .Y(n11925) );
  MUX2X1 U12610 ( .B(ram[2541]), .A(ram[2557]), .S(n12654), .Y(n11895) );
  MUX2X1 U12611 ( .B(ram[2509]), .A(ram[2525]), .S(n12654), .Y(n11894) );
  MUX2X1 U12612 ( .B(ram[2477]), .A(ram[2493]), .S(n12654), .Y(n11898) );
  MUX2X1 U12613 ( .B(ram[2445]), .A(ram[2461]), .S(n12654), .Y(n11897) );
  MUX2X1 U12614 ( .B(n11896), .A(n11893), .S(n12579), .Y(n11907) );
  MUX2X1 U12615 ( .B(ram[2413]), .A(ram[2429]), .S(n12654), .Y(n11901) );
  MUX2X1 U12616 ( .B(ram[2381]), .A(ram[2397]), .S(n12654), .Y(n11900) );
  MUX2X1 U12617 ( .B(ram[2349]), .A(ram[2365]), .S(n12654), .Y(n11904) );
  MUX2X1 U12618 ( .B(ram[2317]), .A(ram[2333]), .S(n12654), .Y(n11903) );
  MUX2X1 U12619 ( .B(n11902), .A(n11899), .S(n12579), .Y(n11906) );
  MUX2X1 U12620 ( .B(ram[2285]), .A(ram[2301]), .S(n12654), .Y(n11910) );
  MUX2X1 U12621 ( .B(ram[2253]), .A(ram[2269]), .S(n12654), .Y(n11909) );
  MUX2X1 U12622 ( .B(ram[2221]), .A(ram[2237]), .S(n12654), .Y(n11913) );
  MUX2X1 U12623 ( .B(ram[2189]), .A(ram[2205]), .S(n12654), .Y(n11912) );
  MUX2X1 U12624 ( .B(n11911), .A(n11908), .S(n12579), .Y(n11922) );
  MUX2X1 U12625 ( .B(ram[2157]), .A(ram[2173]), .S(n12655), .Y(n11916) );
  MUX2X1 U12626 ( .B(ram[2125]), .A(ram[2141]), .S(n12655), .Y(n11915) );
  MUX2X1 U12627 ( .B(ram[2093]), .A(ram[2109]), .S(n12655), .Y(n11919) );
  MUX2X1 U12628 ( .B(ram[2061]), .A(ram[2077]), .S(n12655), .Y(n11918) );
  MUX2X1 U12629 ( .B(n11917), .A(n11914), .S(n12579), .Y(n11921) );
  MUX2X1 U12630 ( .B(n11920), .A(n11905), .S(n12566), .Y(n11924) );
  MUX2X1 U12631 ( .B(n11923), .A(n11860), .S(mem_access_addr[6]), .Y(n12053)
         );
  MUX2X1 U12632 ( .B(ram[2029]), .A(ram[2045]), .S(n12655), .Y(n11928) );
  MUX2X1 U12633 ( .B(ram[1997]), .A(ram[2013]), .S(n12655), .Y(n11927) );
  MUX2X1 U12634 ( .B(ram[1965]), .A(ram[1981]), .S(n12655), .Y(n11931) );
  MUX2X1 U12635 ( .B(ram[1933]), .A(ram[1949]), .S(n12655), .Y(n11930) );
  MUX2X1 U12636 ( .B(n11929), .A(n11926), .S(n12579), .Y(n11940) );
  MUX2X1 U12637 ( .B(ram[1901]), .A(ram[1917]), .S(n12655), .Y(n11934) );
  MUX2X1 U12638 ( .B(ram[1869]), .A(ram[1885]), .S(n12655), .Y(n11933) );
  MUX2X1 U12639 ( .B(ram[1837]), .A(ram[1853]), .S(n12655), .Y(n11937) );
  MUX2X1 U12640 ( .B(ram[1805]), .A(ram[1821]), .S(n12655), .Y(n11936) );
  MUX2X1 U12641 ( .B(n11935), .A(n11932), .S(n12579), .Y(n11939) );
  MUX2X1 U12642 ( .B(ram[1773]), .A(ram[1789]), .S(n12656), .Y(n11943) );
  MUX2X1 U12643 ( .B(ram[1741]), .A(ram[1757]), .S(n12656), .Y(n11942) );
  MUX2X1 U12644 ( .B(ram[1709]), .A(ram[1725]), .S(n12656), .Y(n11946) );
  MUX2X1 U12645 ( .B(ram[1677]), .A(ram[1693]), .S(n12656), .Y(n11945) );
  MUX2X1 U12646 ( .B(n11944), .A(n11941), .S(n12579), .Y(n11955) );
  MUX2X1 U12647 ( .B(ram[1645]), .A(ram[1661]), .S(n12656), .Y(n11949) );
  MUX2X1 U12648 ( .B(ram[1613]), .A(ram[1629]), .S(n12656), .Y(n11948) );
  MUX2X1 U12649 ( .B(ram[1581]), .A(ram[1597]), .S(n12656), .Y(n11952) );
  MUX2X1 U12650 ( .B(ram[1549]), .A(ram[1565]), .S(n12656), .Y(n11951) );
  MUX2X1 U12651 ( .B(n11950), .A(n11947), .S(n12579), .Y(n11954) );
  MUX2X1 U12652 ( .B(n11953), .A(n11938), .S(n12566), .Y(n11988) );
  MUX2X1 U12653 ( .B(ram[1517]), .A(ram[1533]), .S(n12656), .Y(n11958) );
  MUX2X1 U12654 ( .B(ram[1485]), .A(ram[1501]), .S(n12656), .Y(n11957) );
  MUX2X1 U12655 ( .B(ram[1453]), .A(ram[1469]), .S(n12656), .Y(n11961) );
  MUX2X1 U12656 ( .B(ram[1421]), .A(ram[1437]), .S(n12656), .Y(n11960) );
  MUX2X1 U12657 ( .B(n11959), .A(n11956), .S(n12579), .Y(n11970) );
  MUX2X1 U12658 ( .B(ram[1389]), .A(ram[1405]), .S(n12657), .Y(n11964) );
  MUX2X1 U12659 ( .B(ram[1357]), .A(ram[1373]), .S(n12657), .Y(n11963) );
  MUX2X1 U12660 ( .B(ram[1325]), .A(ram[1341]), .S(n12657), .Y(n11967) );
  MUX2X1 U12661 ( .B(ram[1293]), .A(ram[1309]), .S(n12657), .Y(n11966) );
  MUX2X1 U12662 ( .B(n11965), .A(n11962), .S(n12579), .Y(n11969) );
  MUX2X1 U12663 ( .B(ram[1261]), .A(ram[1277]), .S(n12657), .Y(n11973) );
  MUX2X1 U12664 ( .B(ram[1229]), .A(ram[1245]), .S(n12657), .Y(n11972) );
  MUX2X1 U12665 ( .B(ram[1197]), .A(ram[1213]), .S(n12657), .Y(n11976) );
  MUX2X1 U12666 ( .B(ram[1165]), .A(ram[1181]), .S(n12657), .Y(n11975) );
  MUX2X1 U12667 ( .B(n11974), .A(n11971), .S(n12579), .Y(n11985) );
  MUX2X1 U12668 ( .B(ram[1133]), .A(ram[1149]), .S(n12657), .Y(n11979) );
  MUX2X1 U12669 ( .B(ram[1101]), .A(ram[1117]), .S(n12657), .Y(n11978) );
  MUX2X1 U12670 ( .B(ram[1069]), .A(ram[1085]), .S(n12657), .Y(n11982) );
  MUX2X1 U12671 ( .B(ram[1037]), .A(ram[1053]), .S(n12657), .Y(n11981) );
  MUX2X1 U12672 ( .B(n11980), .A(n11977), .S(n12579), .Y(n11984) );
  MUX2X1 U12673 ( .B(n11983), .A(n11968), .S(n12566), .Y(n11987) );
  MUX2X1 U12674 ( .B(ram[1005]), .A(ram[1021]), .S(n12658), .Y(n11991) );
  MUX2X1 U12675 ( .B(ram[973]), .A(ram[989]), .S(n12658), .Y(n11990) );
  MUX2X1 U12676 ( .B(ram[941]), .A(ram[957]), .S(n12658), .Y(n11994) );
  MUX2X1 U12677 ( .B(ram[909]), .A(ram[925]), .S(n12658), .Y(n11993) );
  MUX2X1 U12678 ( .B(n11992), .A(n11989), .S(n12580), .Y(n12003) );
  MUX2X1 U12679 ( .B(ram[877]), .A(ram[893]), .S(n12658), .Y(n11997) );
  MUX2X1 U12680 ( .B(ram[845]), .A(ram[861]), .S(n12658), .Y(n11996) );
  MUX2X1 U12681 ( .B(ram[813]), .A(ram[829]), .S(n12658), .Y(n12000) );
  MUX2X1 U12682 ( .B(ram[781]), .A(ram[797]), .S(n12658), .Y(n11999) );
  MUX2X1 U12683 ( .B(n11998), .A(n11995), .S(n12580), .Y(n12002) );
  MUX2X1 U12684 ( .B(ram[749]), .A(ram[765]), .S(n12658), .Y(n12006) );
  MUX2X1 U12685 ( .B(ram[717]), .A(ram[733]), .S(n12658), .Y(n12005) );
  MUX2X1 U12686 ( .B(ram[685]), .A(ram[701]), .S(n12658), .Y(n12009) );
  MUX2X1 U12687 ( .B(ram[653]), .A(ram[669]), .S(n12658), .Y(n12008) );
  MUX2X1 U12688 ( .B(n12007), .A(n12004), .S(n12580), .Y(n12018) );
  MUX2X1 U12689 ( .B(ram[621]), .A(ram[637]), .S(n12659), .Y(n12012) );
  MUX2X1 U12690 ( .B(ram[589]), .A(ram[605]), .S(n12659), .Y(n12011) );
  MUX2X1 U12691 ( .B(ram[557]), .A(ram[573]), .S(n12659), .Y(n12015) );
  MUX2X1 U12692 ( .B(ram[525]), .A(ram[541]), .S(n12659), .Y(n12014) );
  MUX2X1 U12693 ( .B(n12013), .A(n12010), .S(n12580), .Y(n12017) );
  MUX2X1 U12694 ( .B(n12016), .A(n12001), .S(n12566), .Y(n12051) );
  MUX2X1 U12695 ( .B(ram[493]), .A(ram[509]), .S(n12659), .Y(n12021) );
  MUX2X1 U12696 ( .B(ram[461]), .A(ram[477]), .S(n12659), .Y(n12020) );
  MUX2X1 U12697 ( .B(ram[429]), .A(ram[445]), .S(n12659), .Y(n12024) );
  MUX2X1 U12698 ( .B(ram[397]), .A(ram[413]), .S(n12659), .Y(n12023) );
  MUX2X1 U12699 ( .B(n12022), .A(n12019), .S(n12580), .Y(n12033) );
  MUX2X1 U12700 ( .B(ram[365]), .A(ram[381]), .S(n12659), .Y(n12027) );
  MUX2X1 U12701 ( .B(ram[333]), .A(ram[349]), .S(n12659), .Y(n12026) );
  MUX2X1 U12702 ( .B(ram[301]), .A(ram[317]), .S(n12659), .Y(n12030) );
  MUX2X1 U12703 ( .B(ram[269]), .A(ram[285]), .S(n12659), .Y(n12029) );
  MUX2X1 U12704 ( .B(n12028), .A(n12025), .S(n12580), .Y(n12032) );
  MUX2X1 U12705 ( .B(ram[237]), .A(ram[253]), .S(n12660), .Y(n12036) );
  MUX2X1 U12706 ( .B(ram[205]), .A(ram[221]), .S(n12660), .Y(n12035) );
  MUX2X1 U12707 ( .B(ram[173]), .A(ram[189]), .S(n12660), .Y(n12039) );
  MUX2X1 U12708 ( .B(ram[141]), .A(ram[157]), .S(n12660), .Y(n12038) );
  MUX2X1 U12709 ( .B(n12037), .A(n12034), .S(n12580), .Y(n12048) );
  MUX2X1 U12710 ( .B(ram[109]), .A(ram[125]), .S(n12660), .Y(n12042) );
  MUX2X1 U12711 ( .B(ram[77]), .A(ram[93]), .S(n12660), .Y(n12041) );
  MUX2X1 U12712 ( .B(ram[45]), .A(ram[61]), .S(n12660), .Y(n12045) );
  MUX2X1 U12713 ( .B(ram[13]), .A(ram[29]), .S(n12660), .Y(n12044) );
  MUX2X1 U12714 ( .B(n12043), .A(n12040), .S(n12580), .Y(n12047) );
  MUX2X1 U12715 ( .B(n12046), .A(n12031), .S(n12566), .Y(n12050) );
  MUX2X1 U12716 ( .B(n12049), .A(n11986), .S(mem_access_addr[6]), .Y(n12052)
         );
  MUX2X1 U12717 ( .B(ram[4078]), .A(ram[4094]), .S(n12660), .Y(n12056) );
  MUX2X1 U12718 ( .B(ram[4046]), .A(ram[4062]), .S(n12660), .Y(n12055) );
  MUX2X1 U12719 ( .B(ram[4014]), .A(ram[4030]), .S(n12660), .Y(n12059) );
  MUX2X1 U12720 ( .B(ram[3982]), .A(ram[3998]), .S(n12660), .Y(n12058) );
  MUX2X1 U12721 ( .B(n12057), .A(n12054), .S(n12580), .Y(n12068) );
  MUX2X1 U12722 ( .B(ram[3950]), .A(ram[3966]), .S(n12661), .Y(n12062) );
  MUX2X1 U12723 ( .B(ram[3918]), .A(ram[3934]), .S(n12661), .Y(n12061) );
  MUX2X1 U12724 ( .B(ram[3886]), .A(ram[3902]), .S(n12661), .Y(n12065) );
  MUX2X1 U12725 ( .B(ram[3854]), .A(ram[3870]), .S(n12661), .Y(n12064) );
  MUX2X1 U12726 ( .B(n12063), .A(n12060), .S(n12580), .Y(n12067) );
  MUX2X1 U12727 ( .B(ram[3822]), .A(ram[3838]), .S(n12661), .Y(n12071) );
  MUX2X1 U12728 ( .B(ram[3790]), .A(ram[3806]), .S(n12661), .Y(n12070) );
  MUX2X1 U12729 ( .B(ram[3758]), .A(ram[3774]), .S(n12661), .Y(n12074) );
  MUX2X1 U12730 ( .B(ram[3726]), .A(ram[3742]), .S(n12661), .Y(n12073) );
  MUX2X1 U12731 ( .B(n12072), .A(n12069), .S(n12580), .Y(n12083) );
  MUX2X1 U12732 ( .B(ram[3694]), .A(ram[3710]), .S(n12661), .Y(n12077) );
  MUX2X1 U12733 ( .B(ram[3662]), .A(ram[3678]), .S(n12661), .Y(n12076) );
  MUX2X1 U12734 ( .B(ram[3630]), .A(ram[3646]), .S(n12661), .Y(n12080) );
  MUX2X1 U12735 ( .B(ram[3598]), .A(ram[3614]), .S(n12661), .Y(n12079) );
  MUX2X1 U12736 ( .B(n12078), .A(n12075), .S(n12580), .Y(n12082) );
  MUX2X1 U12737 ( .B(n12081), .A(n12066), .S(n12566), .Y(n12116) );
  MUX2X1 U12738 ( .B(ram[3566]), .A(ram[3582]), .S(n12662), .Y(n12086) );
  MUX2X1 U12739 ( .B(ram[3534]), .A(ram[3550]), .S(n12662), .Y(n12085) );
  MUX2X1 U12740 ( .B(ram[3502]), .A(ram[3518]), .S(n12662), .Y(n12089) );
  MUX2X1 U12741 ( .B(ram[3470]), .A(ram[3486]), .S(n12662), .Y(n12088) );
  MUX2X1 U12742 ( .B(n12087), .A(n12084), .S(n12581), .Y(n12098) );
  MUX2X1 U12743 ( .B(ram[3438]), .A(ram[3454]), .S(n12662), .Y(n12092) );
  MUX2X1 U12744 ( .B(ram[3406]), .A(ram[3422]), .S(n12662), .Y(n12091) );
  MUX2X1 U12745 ( .B(ram[3374]), .A(ram[3390]), .S(n12662), .Y(n12095) );
  MUX2X1 U12746 ( .B(ram[3342]), .A(ram[3358]), .S(n12662), .Y(n12094) );
  MUX2X1 U12747 ( .B(n12093), .A(n12090), .S(n12581), .Y(n12097) );
  MUX2X1 U12748 ( .B(ram[3310]), .A(ram[3326]), .S(n12662), .Y(n12101) );
  MUX2X1 U12749 ( .B(ram[3278]), .A(ram[3294]), .S(n12662), .Y(n12100) );
  MUX2X1 U12750 ( .B(ram[3246]), .A(ram[3262]), .S(n12662), .Y(n12104) );
  MUX2X1 U12751 ( .B(ram[3214]), .A(ram[3230]), .S(n12662), .Y(n12103) );
  MUX2X1 U12752 ( .B(n12102), .A(n12099), .S(n12581), .Y(n12113) );
  MUX2X1 U12753 ( .B(ram[3182]), .A(ram[3198]), .S(n12663), .Y(n12107) );
  MUX2X1 U12754 ( .B(ram[3150]), .A(ram[3166]), .S(n12663), .Y(n12106) );
  MUX2X1 U12755 ( .B(ram[3118]), .A(ram[3134]), .S(n12663), .Y(n12110) );
  MUX2X1 U12756 ( .B(ram[3086]), .A(ram[3102]), .S(n12663), .Y(n12109) );
  MUX2X1 U12757 ( .B(n12108), .A(n12105), .S(n12581), .Y(n12112) );
  MUX2X1 U12758 ( .B(n12111), .A(n12096), .S(n12566), .Y(n12115) );
  MUX2X1 U12759 ( .B(ram[3054]), .A(ram[3070]), .S(n12663), .Y(n12119) );
  MUX2X1 U12760 ( .B(ram[3022]), .A(ram[3038]), .S(n12663), .Y(n12118) );
  MUX2X1 U12761 ( .B(ram[2990]), .A(ram[3006]), .S(n12663), .Y(n12122) );
  MUX2X1 U12762 ( .B(ram[2958]), .A(ram[2974]), .S(n12663), .Y(n12121) );
  MUX2X1 U12763 ( .B(n12120), .A(n12117), .S(n12581), .Y(n12131) );
  MUX2X1 U12764 ( .B(ram[2926]), .A(ram[2942]), .S(n12663), .Y(n12125) );
  MUX2X1 U12765 ( .B(ram[2894]), .A(ram[2910]), .S(n12663), .Y(n12124) );
  MUX2X1 U12766 ( .B(ram[2862]), .A(ram[2878]), .S(n12663), .Y(n12128) );
  MUX2X1 U12767 ( .B(ram[2830]), .A(ram[2846]), .S(n12663), .Y(n12127) );
  MUX2X1 U12768 ( .B(n12126), .A(n12123), .S(n12581), .Y(n12130) );
  MUX2X1 U12769 ( .B(ram[2798]), .A(ram[2814]), .S(n12664), .Y(n12134) );
  MUX2X1 U12770 ( .B(ram[2766]), .A(ram[2782]), .S(n12664), .Y(n12133) );
  MUX2X1 U12771 ( .B(ram[2734]), .A(ram[2750]), .S(n12664), .Y(n12137) );
  MUX2X1 U12772 ( .B(ram[2702]), .A(ram[2718]), .S(n12664), .Y(n12136) );
  MUX2X1 U12773 ( .B(n12135), .A(n12132), .S(n12581), .Y(n12146) );
  MUX2X1 U12774 ( .B(ram[2670]), .A(ram[2686]), .S(n12664), .Y(n12140) );
  MUX2X1 U12775 ( .B(ram[2638]), .A(ram[2654]), .S(n12664), .Y(n12139) );
  MUX2X1 U12776 ( .B(ram[2606]), .A(ram[2622]), .S(n12664), .Y(n12143) );
  MUX2X1 U12777 ( .B(ram[2574]), .A(ram[2590]), .S(n12664), .Y(n12142) );
  MUX2X1 U12778 ( .B(n12141), .A(n12138), .S(n12581), .Y(n12145) );
  MUX2X1 U12779 ( .B(n12144), .A(n12129), .S(n12566), .Y(n12179) );
  MUX2X1 U12780 ( .B(ram[2542]), .A(ram[2558]), .S(n12664), .Y(n12149) );
  MUX2X1 U12781 ( .B(ram[2510]), .A(ram[2526]), .S(n12664), .Y(n12148) );
  MUX2X1 U12782 ( .B(ram[2478]), .A(ram[2494]), .S(n12664), .Y(n12152) );
  MUX2X1 U12783 ( .B(ram[2446]), .A(ram[2462]), .S(n12664), .Y(n12151) );
  MUX2X1 U12784 ( .B(n12150), .A(n12147), .S(n12581), .Y(n12161) );
  MUX2X1 U12785 ( .B(ram[2414]), .A(ram[2430]), .S(n12665), .Y(n12155) );
  MUX2X1 U12786 ( .B(ram[2382]), .A(ram[2398]), .S(n12665), .Y(n12154) );
  MUX2X1 U12787 ( .B(ram[2350]), .A(ram[2366]), .S(n12665), .Y(n12158) );
  MUX2X1 U12788 ( .B(ram[2318]), .A(ram[2334]), .S(n12665), .Y(n12157) );
  MUX2X1 U12789 ( .B(n12156), .A(n12153), .S(n12581), .Y(n12160) );
  MUX2X1 U12790 ( .B(ram[2286]), .A(ram[2302]), .S(n12665), .Y(n12164) );
  MUX2X1 U12791 ( .B(ram[2254]), .A(ram[2270]), .S(n12665), .Y(n12163) );
  MUX2X1 U12792 ( .B(ram[2222]), .A(ram[2238]), .S(n12665), .Y(n12167) );
  MUX2X1 U12793 ( .B(ram[2190]), .A(ram[2206]), .S(n12665), .Y(n12166) );
  MUX2X1 U12794 ( .B(n12165), .A(n12162), .S(n12581), .Y(n12176) );
  MUX2X1 U12795 ( .B(ram[2158]), .A(ram[2174]), .S(n12665), .Y(n12170) );
  MUX2X1 U12796 ( .B(ram[2126]), .A(ram[2142]), .S(n12665), .Y(n12169) );
  MUX2X1 U12797 ( .B(ram[2094]), .A(ram[2110]), .S(n12665), .Y(n12173) );
  MUX2X1 U12798 ( .B(ram[2062]), .A(ram[2078]), .S(n12665), .Y(n12172) );
  MUX2X1 U12799 ( .B(n12171), .A(n12168), .S(n12581), .Y(n12175) );
  MUX2X1 U12800 ( .B(n12174), .A(n12159), .S(n12566), .Y(n12178) );
  MUX2X1 U12801 ( .B(n12177), .A(n12114), .S(mem_access_addr[6]), .Y(n12307)
         );
  MUX2X1 U12802 ( .B(ram[2030]), .A(ram[2046]), .S(n12666), .Y(n12182) );
  MUX2X1 U12803 ( .B(ram[1998]), .A(ram[2014]), .S(n12666), .Y(n12181) );
  MUX2X1 U12804 ( .B(ram[1966]), .A(ram[1982]), .S(n12666), .Y(n12185) );
  MUX2X1 U12805 ( .B(ram[1934]), .A(ram[1950]), .S(n12666), .Y(n12184) );
  MUX2X1 U12806 ( .B(n12183), .A(n12180), .S(n12582), .Y(n12194) );
  MUX2X1 U12807 ( .B(ram[1902]), .A(ram[1918]), .S(n12666), .Y(n12188) );
  MUX2X1 U12808 ( .B(ram[1870]), .A(ram[1886]), .S(n12666), .Y(n12187) );
  MUX2X1 U12809 ( .B(ram[1838]), .A(ram[1854]), .S(n12666), .Y(n12191) );
  MUX2X1 U12810 ( .B(ram[1806]), .A(ram[1822]), .S(n12666), .Y(n12190) );
  MUX2X1 U12811 ( .B(n12189), .A(n12186), .S(n12582), .Y(n12193) );
  MUX2X1 U12812 ( .B(ram[1774]), .A(ram[1790]), .S(n12666), .Y(n12197) );
  MUX2X1 U12813 ( .B(ram[1742]), .A(ram[1758]), .S(n12666), .Y(n12196) );
  MUX2X1 U12814 ( .B(ram[1710]), .A(ram[1726]), .S(n12666), .Y(n12200) );
  MUX2X1 U12815 ( .B(ram[1678]), .A(ram[1694]), .S(n12666), .Y(n12199) );
  MUX2X1 U12816 ( .B(n12198), .A(n12195), .S(n12582), .Y(n12209) );
  MUX2X1 U12817 ( .B(ram[1646]), .A(ram[1662]), .S(n12667), .Y(n12203) );
  MUX2X1 U12818 ( .B(ram[1614]), .A(ram[1630]), .S(n12667), .Y(n12202) );
  MUX2X1 U12819 ( .B(ram[1582]), .A(ram[1598]), .S(n12667), .Y(n12206) );
  MUX2X1 U12820 ( .B(ram[1550]), .A(ram[1566]), .S(n12667), .Y(n12205) );
  MUX2X1 U12821 ( .B(n12204), .A(n12201), .S(n12582), .Y(n12208) );
  MUX2X1 U12822 ( .B(n12207), .A(n12192), .S(n12567), .Y(n12242) );
  MUX2X1 U12823 ( .B(ram[1518]), .A(ram[1534]), .S(n12667), .Y(n12212) );
  MUX2X1 U12824 ( .B(ram[1486]), .A(ram[1502]), .S(n12667), .Y(n12211) );
  MUX2X1 U12825 ( .B(ram[1454]), .A(ram[1470]), .S(n12667), .Y(n12215) );
  MUX2X1 U12826 ( .B(ram[1422]), .A(ram[1438]), .S(n12667), .Y(n12214) );
  MUX2X1 U12827 ( .B(n12213), .A(n12210), .S(n12582), .Y(n12224) );
  MUX2X1 U12828 ( .B(ram[1390]), .A(ram[1406]), .S(n12667), .Y(n12218) );
  MUX2X1 U12829 ( .B(ram[1358]), .A(ram[1374]), .S(n12667), .Y(n12217) );
  MUX2X1 U12830 ( .B(ram[1326]), .A(ram[1342]), .S(n12667), .Y(n12221) );
  MUX2X1 U12831 ( .B(ram[1294]), .A(ram[1310]), .S(n12667), .Y(n12220) );
  MUX2X1 U12832 ( .B(n12219), .A(n12216), .S(n12582), .Y(n12223) );
  MUX2X1 U12833 ( .B(ram[1262]), .A(ram[1278]), .S(n12668), .Y(n12227) );
  MUX2X1 U12834 ( .B(ram[1230]), .A(ram[1246]), .S(n12668), .Y(n12226) );
  MUX2X1 U12835 ( .B(ram[1198]), .A(ram[1214]), .S(n12668), .Y(n12230) );
  MUX2X1 U12836 ( .B(ram[1166]), .A(ram[1182]), .S(n12668), .Y(n12229) );
  MUX2X1 U12837 ( .B(n12228), .A(n12225), .S(n12582), .Y(n12239) );
  MUX2X1 U12838 ( .B(ram[1134]), .A(ram[1150]), .S(n12668), .Y(n12233) );
  MUX2X1 U12839 ( .B(ram[1102]), .A(ram[1118]), .S(n12668), .Y(n12232) );
  MUX2X1 U12840 ( .B(ram[1070]), .A(ram[1086]), .S(n12668), .Y(n12236) );
  MUX2X1 U12841 ( .B(ram[1038]), .A(ram[1054]), .S(n12668), .Y(n12235) );
  MUX2X1 U12842 ( .B(n12234), .A(n12231), .S(n12582), .Y(n12238) );
  MUX2X1 U12843 ( .B(n12237), .A(n12222), .S(n12567), .Y(n12241) );
  MUX2X1 U12844 ( .B(ram[1006]), .A(ram[1022]), .S(n12668), .Y(n12245) );
  MUX2X1 U12845 ( .B(ram[974]), .A(ram[990]), .S(n12668), .Y(n12244) );
  MUX2X1 U12846 ( .B(ram[942]), .A(ram[958]), .S(n12668), .Y(n12248) );
  MUX2X1 U12847 ( .B(ram[910]), .A(ram[926]), .S(n12668), .Y(n12247) );
  MUX2X1 U12848 ( .B(n12246), .A(n12243), .S(n12582), .Y(n12257) );
  MUX2X1 U12849 ( .B(ram[878]), .A(ram[894]), .S(n12669), .Y(n12251) );
  MUX2X1 U12850 ( .B(ram[846]), .A(ram[862]), .S(n12669), .Y(n12250) );
  MUX2X1 U12851 ( .B(ram[814]), .A(ram[830]), .S(n12669), .Y(n12254) );
  MUX2X1 U12852 ( .B(ram[782]), .A(ram[798]), .S(n12669), .Y(n12253) );
  MUX2X1 U12853 ( .B(n12252), .A(n12249), .S(n12582), .Y(n12256) );
  MUX2X1 U12854 ( .B(ram[750]), .A(ram[766]), .S(n12669), .Y(n12260) );
  MUX2X1 U12855 ( .B(ram[718]), .A(ram[734]), .S(n12669), .Y(n12259) );
  MUX2X1 U12856 ( .B(ram[686]), .A(ram[702]), .S(n12669), .Y(n12263) );
  MUX2X1 U12857 ( .B(ram[654]), .A(ram[670]), .S(n12669), .Y(n12262) );
  MUX2X1 U12858 ( .B(n12261), .A(n12258), .S(n12582), .Y(n12272) );
  MUX2X1 U12859 ( .B(ram[622]), .A(ram[638]), .S(n12669), .Y(n12266) );
  MUX2X1 U12860 ( .B(ram[590]), .A(ram[606]), .S(n12669), .Y(n12265) );
  MUX2X1 U12861 ( .B(ram[558]), .A(ram[574]), .S(n12669), .Y(n12269) );
  MUX2X1 U12862 ( .B(ram[526]), .A(ram[542]), .S(n12669), .Y(n12268) );
  MUX2X1 U12863 ( .B(n12267), .A(n12264), .S(n12582), .Y(n12271) );
  MUX2X1 U12864 ( .B(n12270), .A(n12255), .S(n12567), .Y(n12305) );
  MUX2X1 U12865 ( .B(ram[494]), .A(ram[510]), .S(n12670), .Y(n12275) );
  MUX2X1 U12866 ( .B(ram[462]), .A(ram[478]), .S(n12670), .Y(n12274) );
  MUX2X1 U12867 ( .B(ram[430]), .A(ram[446]), .S(n12670), .Y(n12278) );
  MUX2X1 U12868 ( .B(ram[398]), .A(ram[414]), .S(n12670), .Y(n12277) );
  MUX2X1 U12869 ( .B(n12276), .A(n12273), .S(n12583), .Y(n12287) );
  MUX2X1 U12870 ( .B(ram[366]), .A(ram[382]), .S(n12670), .Y(n12281) );
  MUX2X1 U12871 ( .B(ram[334]), .A(ram[350]), .S(n12670), .Y(n12280) );
  MUX2X1 U12872 ( .B(ram[302]), .A(ram[318]), .S(n12670), .Y(n12284) );
  MUX2X1 U12873 ( .B(ram[270]), .A(ram[286]), .S(n12670), .Y(n12283) );
  MUX2X1 U12874 ( .B(n12282), .A(n12279), .S(n12583), .Y(n12286) );
  MUX2X1 U12875 ( .B(ram[238]), .A(ram[254]), .S(n12670), .Y(n12290) );
  MUX2X1 U12876 ( .B(ram[206]), .A(ram[222]), .S(n12670), .Y(n12289) );
  MUX2X1 U12877 ( .B(ram[174]), .A(ram[190]), .S(n12670), .Y(n12293) );
  MUX2X1 U12878 ( .B(ram[142]), .A(ram[158]), .S(n12670), .Y(n12292) );
  MUX2X1 U12879 ( .B(n12291), .A(n12288), .S(n12583), .Y(n12302) );
  MUX2X1 U12880 ( .B(ram[110]), .A(ram[126]), .S(n12671), .Y(n12296) );
  MUX2X1 U12881 ( .B(ram[78]), .A(ram[94]), .S(n12671), .Y(n12295) );
  MUX2X1 U12882 ( .B(ram[46]), .A(ram[62]), .S(n12671), .Y(n12299) );
  MUX2X1 U12883 ( .B(ram[14]), .A(ram[30]), .S(n12671), .Y(n12298) );
  MUX2X1 U12884 ( .B(n12297), .A(n12294), .S(n12583), .Y(n12301) );
  MUX2X1 U12885 ( .B(n12300), .A(n12285), .S(n12567), .Y(n12304) );
  MUX2X1 U12886 ( .B(n12303), .A(n12240), .S(mem_access_addr[6]), .Y(n12306)
         );
  MUX2X1 U12887 ( .B(ram[4079]), .A(ram[4095]), .S(n12671), .Y(n12310) );
  MUX2X1 U12888 ( .B(ram[4047]), .A(ram[4063]), .S(n12671), .Y(n12309) );
  MUX2X1 U12889 ( .B(ram[4015]), .A(ram[4031]), .S(n12671), .Y(n12313) );
  MUX2X1 U12890 ( .B(ram[3983]), .A(ram[3999]), .S(n12671), .Y(n12312) );
  MUX2X1 U12891 ( .B(n12311), .A(n12308), .S(n12583), .Y(n12322) );
  MUX2X1 U12892 ( .B(ram[3951]), .A(ram[3967]), .S(n12671), .Y(n12316) );
  MUX2X1 U12893 ( .B(ram[3919]), .A(ram[3935]), .S(n12671), .Y(n12315) );
  MUX2X1 U12894 ( .B(ram[3887]), .A(ram[3903]), .S(n12671), .Y(n12319) );
  MUX2X1 U12895 ( .B(ram[3855]), .A(ram[3871]), .S(n12671), .Y(n12318) );
  MUX2X1 U12896 ( .B(n12317), .A(n12314), .S(n12583), .Y(n12321) );
  MUX2X1 U12897 ( .B(ram[3823]), .A(ram[3839]), .S(n12672), .Y(n12325) );
  MUX2X1 U12898 ( .B(ram[3791]), .A(ram[3807]), .S(n12672), .Y(n12324) );
  MUX2X1 U12899 ( .B(ram[3759]), .A(ram[3775]), .S(n12672), .Y(n12328) );
  MUX2X1 U12900 ( .B(ram[3727]), .A(ram[3743]), .S(n12672), .Y(n12327) );
  MUX2X1 U12901 ( .B(n12326), .A(n12323), .S(n12583), .Y(n12337) );
  MUX2X1 U12902 ( .B(ram[3695]), .A(ram[3711]), .S(n12672), .Y(n12331) );
  MUX2X1 U12903 ( .B(ram[3663]), .A(ram[3679]), .S(n12672), .Y(n12330) );
  MUX2X1 U12904 ( .B(ram[3631]), .A(ram[3647]), .S(n12672), .Y(n12334) );
  MUX2X1 U12905 ( .B(ram[3599]), .A(ram[3615]), .S(n12672), .Y(n12333) );
  MUX2X1 U12906 ( .B(n12332), .A(n12329), .S(n12583), .Y(n12336) );
  MUX2X1 U12907 ( .B(n12335), .A(n12320), .S(n12567), .Y(n12370) );
  MUX2X1 U12908 ( .B(ram[3567]), .A(ram[3583]), .S(n12672), .Y(n12340) );
  MUX2X1 U12909 ( .B(ram[3535]), .A(ram[3551]), .S(n12672), .Y(n12339) );
  MUX2X1 U12910 ( .B(ram[3503]), .A(ram[3519]), .S(n12672), .Y(n12343) );
  MUX2X1 U12911 ( .B(ram[3471]), .A(ram[3487]), .S(n12672), .Y(n12342) );
  MUX2X1 U12912 ( .B(n12341), .A(n12338), .S(n12583), .Y(n12352) );
  MUX2X1 U12913 ( .B(ram[3439]), .A(ram[3455]), .S(n12673), .Y(n12346) );
  MUX2X1 U12914 ( .B(ram[3407]), .A(ram[3423]), .S(n12673), .Y(n12345) );
  MUX2X1 U12915 ( .B(ram[3375]), .A(ram[3391]), .S(n12673), .Y(n12349) );
  MUX2X1 U12916 ( .B(ram[3343]), .A(ram[3359]), .S(n12673), .Y(n12348) );
  MUX2X1 U12917 ( .B(n12347), .A(n12344), .S(n12583), .Y(n12351) );
  MUX2X1 U12918 ( .B(ram[3311]), .A(ram[3327]), .S(n12673), .Y(n12355) );
  MUX2X1 U12919 ( .B(ram[3279]), .A(ram[3295]), .S(n12673), .Y(n12354) );
  MUX2X1 U12920 ( .B(ram[3247]), .A(ram[3263]), .S(n12673), .Y(n12358) );
  MUX2X1 U12921 ( .B(ram[3215]), .A(ram[3231]), .S(n12673), .Y(n12357) );
  MUX2X1 U12922 ( .B(n12356), .A(n12353), .S(n12583), .Y(n12367) );
  MUX2X1 U12923 ( .B(ram[3183]), .A(ram[3199]), .S(n12673), .Y(n12361) );
  MUX2X1 U12924 ( .B(ram[3151]), .A(ram[3167]), .S(n12673), .Y(n12360) );
  MUX2X1 U12925 ( .B(ram[3119]), .A(ram[3135]), .S(n12673), .Y(n12364) );
  MUX2X1 U12926 ( .B(ram[3087]), .A(ram[3103]), .S(n12673), .Y(n12363) );
  MUX2X1 U12927 ( .B(n12362), .A(n12359), .S(n12583), .Y(n12366) );
  MUX2X1 U12928 ( .B(n12365), .A(n12350), .S(n12567), .Y(n12369) );
  MUX2X1 U12929 ( .B(ram[3055]), .A(ram[3071]), .S(n12674), .Y(n12373) );
  MUX2X1 U12930 ( .B(ram[3023]), .A(ram[3039]), .S(n12674), .Y(n12372) );
  MUX2X1 U12931 ( .B(ram[2991]), .A(ram[3007]), .S(n12674), .Y(n12376) );
  MUX2X1 U12932 ( .B(ram[2959]), .A(ram[2975]), .S(n12674), .Y(n12375) );
  MUX2X1 U12933 ( .B(n12374), .A(n12371), .S(n12584), .Y(n12385) );
  MUX2X1 U12934 ( .B(ram[2927]), .A(ram[2943]), .S(n12674), .Y(n12379) );
  MUX2X1 U12935 ( .B(ram[2895]), .A(ram[2911]), .S(n12674), .Y(n12378) );
  MUX2X1 U12936 ( .B(ram[2863]), .A(ram[2879]), .S(n12674), .Y(n12382) );
  MUX2X1 U12937 ( .B(ram[2831]), .A(ram[2847]), .S(n12674), .Y(n12381) );
  MUX2X1 U12938 ( .B(n12380), .A(n12377), .S(n12584), .Y(n12384) );
  MUX2X1 U12939 ( .B(ram[2799]), .A(ram[2815]), .S(n12674), .Y(n12388) );
  MUX2X1 U12940 ( .B(ram[2767]), .A(ram[2783]), .S(n12674), .Y(n12387) );
  MUX2X1 U12941 ( .B(ram[2735]), .A(ram[2751]), .S(n12674), .Y(n12391) );
  MUX2X1 U12942 ( .B(ram[2703]), .A(ram[2719]), .S(n12674), .Y(n12390) );
  MUX2X1 U12943 ( .B(n12389), .A(n12386), .S(n12584), .Y(n12400) );
  MUX2X1 U12944 ( .B(ram[2671]), .A(ram[2687]), .S(n12675), .Y(n12394) );
  MUX2X1 U12945 ( .B(ram[2639]), .A(ram[2655]), .S(n12675), .Y(n12393) );
  MUX2X1 U12946 ( .B(ram[2607]), .A(ram[2623]), .S(n12675), .Y(n12397) );
  MUX2X1 U12947 ( .B(ram[2575]), .A(ram[2591]), .S(n12675), .Y(n12396) );
  MUX2X1 U12948 ( .B(n12395), .A(n12392), .S(n12584), .Y(n12399) );
  MUX2X1 U12949 ( .B(n12398), .A(n12383), .S(n12567), .Y(n12433) );
  MUX2X1 U12950 ( .B(ram[2543]), .A(ram[2559]), .S(n12675), .Y(n12403) );
  MUX2X1 U12951 ( .B(ram[2511]), .A(ram[2527]), .S(n12675), .Y(n12402) );
  MUX2X1 U12952 ( .B(ram[2479]), .A(ram[2495]), .S(n12675), .Y(n12406) );
  MUX2X1 U12953 ( .B(ram[2447]), .A(ram[2463]), .S(n12675), .Y(n12405) );
  MUX2X1 U12954 ( .B(n12404), .A(n12401), .S(n12584), .Y(n12415) );
  MUX2X1 U12955 ( .B(ram[2415]), .A(ram[2431]), .S(n12675), .Y(n12409) );
  MUX2X1 U12956 ( .B(ram[2383]), .A(ram[2399]), .S(n12675), .Y(n12408) );
  MUX2X1 U12957 ( .B(ram[2351]), .A(ram[2367]), .S(n12675), .Y(n12412) );
  MUX2X1 U12958 ( .B(ram[2319]), .A(ram[2335]), .S(n12675), .Y(n12411) );
  MUX2X1 U12959 ( .B(n12410), .A(n12407), .S(n12584), .Y(n12414) );
  MUX2X1 U12960 ( .B(ram[2287]), .A(ram[2303]), .S(n12676), .Y(n12418) );
  MUX2X1 U12961 ( .B(ram[2255]), .A(ram[2271]), .S(n12676), .Y(n12417) );
  MUX2X1 U12962 ( .B(ram[2223]), .A(ram[2239]), .S(n12676), .Y(n12421) );
  MUX2X1 U12963 ( .B(ram[2191]), .A(ram[2207]), .S(n12676), .Y(n12420) );
  MUX2X1 U12964 ( .B(n12419), .A(n12416), .S(n12584), .Y(n12430) );
  MUX2X1 U12965 ( .B(ram[2159]), .A(ram[2175]), .S(n12676), .Y(n12424) );
  MUX2X1 U12966 ( .B(ram[2127]), .A(ram[2143]), .S(n12676), .Y(n12423) );
  MUX2X1 U12967 ( .B(ram[2095]), .A(ram[2111]), .S(n12676), .Y(n12427) );
  MUX2X1 U12968 ( .B(ram[2063]), .A(ram[2079]), .S(n12676), .Y(n12426) );
  MUX2X1 U12969 ( .B(n12425), .A(n12422), .S(n12584), .Y(n12429) );
  MUX2X1 U12970 ( .B(n12428), .A(n12413), .S(n12567), .Y(n12432) );
  MUX2X1 U12971 ( .B(n12431), .A(n12368), .S(mem_access_addr[6]), .Y(n12561)
         );
  MUX2X1 U12972 ( .B(ram[2031]), .A(ram[2047]), .S(n12676), .Y(n12436) );
  MUX2X1 U12973 ( .B(ram[1999]), .A(ram[2015]), .S(n12676), .Y(n12435) );
  MUX2X1 U12974 ( .B(ram[1967]), .A(ram[1983]), .S(n12676), .Y(n12439) );
  MUX2X1 U12975 ( .B(ram[1935]), .A(ram[1951]), .S(n12676), .Y(n12438) );
  MUX2X1 U12976 ( .B(n12437), .A(n12434), .S(n12584), .Y(n12448) );
  MUX2X1 U12977 ( .B(ram[1903]), .A(ram[1919]), .S(n12677), .Y(n12442) );
  MUX2X1 U12978 ( .B(ram[1871]), .A(ram[1887]), .S(n12677), .Y(n12441) );
  MUX2X1 U12979 ( .B(ram[1839]), .A(ram[1855]), .S(n12677), .Y(n12445) );
  MUX2X1 U12980 ( .B(ram[1807]), .A(ram[1823]), .S(n12677), .Y(n12444) );
  MUX2X1 U12981 ( .B(n12443), .A(n12440), .S(n12584), .Y(n12447) );
  MUX2X1 U12982 ( .B(ram[1775]), .A(ram[1791]), .S(n12677), .Y(n12451) );
  MUX2X1 U12983 ( .B(ram[1743]), .A(ram[1759]), .S(n12677), .Y(n12450) );
  MUX2X1 U12984 ( .B(ram[1711]), .A(ram[1727]), .S(n12677), .Y(n12454) );
  MUX2X1 U12985 ( .B(ram[1679]), .A(ram[1695]), .S(n12677), .Y(n12453) );
  MUX2X1 U12986 ( .B(n12452), .A(n12449), .S(n12584), .Y(n12463) );
  MUX2X1 U12987 ( .B(ram[1647]), .A(ram[1663]), .S(n12677), .Y(n12457) );
  MUX2X1 U12988 ( .B(ram[1615]), .A(ram[1631]), .S(n12677), .Y(n12456) );
  MUX2X1 U12989 ( .B(ram[1583]), .A(ram[1599]), .S(n12677), .Y(n12460) );
  MUX2X1 U12990 ( .B(ram[1551]), .A(ram[1567]), .S(n12677), .Y(n12459) );
  MUX2X1 U12991 ( .B(n12458), .A(n12455), .S(n12584), .Y(n12462) );
  MUX2X1 U12992 ( .B(n12461), .A(n12446), .S(n12567), .Y(n12496) );
  MUX2X1 U12993 ( .B(ram[1519]), .A(ram[1535]), .S(n12678), .Y(n12466) );
  MUX2X1 U12994 ( .B(ram[1487]), .A(ram[1503]), .S(n12678), .Y(n12465) );
  MUX2X1 U12995 ( .B(ram[1455]), .A(ram[1471]), .S(n12678), .Y(n12469) );
  MUX2X1 U12996 ( .B(ram[1423]), .A(ram[1439]), .S(n12678), .Y(n12468) );
  MUX2X1 U12997 ( .B(n12467), .A(n12464), .S(n12585), .Y(n12478) );
  MUX2X1 U12998 ( .B(ram[1391]), .A(ram[1407]), .S(n12678), .Y(n12472) );
  MUX2X1 U12999 ( .B(ram[1359]), .A(ram[1375]), .S(n12678), .Y(n12471) );
  MUX2X1 U13000 ( .B(ram[1327]), .A(ram[1343]), .S(n12678), .Y(n12475) );
  MUX2X1 U13001 ( .B(ram[1295]), .A(ram[1311]), .S(n12678), .Y(n12474) );
  MUX2X1 U13002 ( .B(n12473), .A(n12470), .S(n12585), .Y(n12477) );
  MUX2X1 U13003 ( .B(ram[1263]), .A(ram[1279]), .S(n12678), .Y(n12481) );
  MUX2X1 U13004 ( .B(ram[1231]), .A(ram[1247]), .S(n12678), .Y(n12480) );
  MUX2X1 U13005 ( .B(ram[1199]), .A(ram[1215]), .S(n12678), .Y(n12484) );
  MUX2X1 U13006 ( .B(ram[1167]), .A(ram[1183]), .S(n12678), .Y(n12483) );
  MUX2X1 U13007 ( .B(n12482), .A(n12479), .S(n12585), .Y(n12493) );
  MUX2X1 U13008 ( .B(ram[1135]), .A(ram[1151]), .S(n12679), .Y(n12487) );
  MUX2X1 U13009 ( .B(ram[1103]), .A(ram[1119]), .S(n12679), .Y(n12486) );
  MUX2X1 U13010 ( .B(ram[1071]), .A(ram[1087]), .S(n12679), .Y(n12490) );
  MUX2X1 U13011 ( .B(ram[1039]), .A(ram[1055]), .S(n12679), .Y(n12489) );
  MUX2X1 U13012 ( .B(n12488), .A(n12485), .S(n12585), .Y(n12492) );
  MUX2X1 U13013 ( .B(n12491), .A(n12476), .S(n12567), .Y(n12495) );
  MUX2X1 U13014 ( .B(ram[1007]), .A(ram[1023]), .S(n12679), .Y(n12499) );
  MUX2X1 U13015 ( .B(ram[975]), .A(ram[991]), .S(n12679), .Y(n12498) );
  MUX2X1 U13016 ( .B(ram[943]), .A(ram[959]), .S(n12679), .Y(n12502) );
  MUX2X1 U13017 ( .B(ram[911]), .A(ram[927]), .S(n12679), .Y(n12501) );
  MUX2X1 U13018 ( .B(n12500), .A(n12497), .S(n12585), .Y(n12511) );
  MUX2X1 U13019 ( .B(ram[879]), .A(ram[895]), .S(n12679), .Y(n12505) );
  MUX2X1 U13020 ( .B(ram[847]), .A(ram[863]), .S(n12679), .Y(n12504) );
  MUX2X1 U13021 ( .B(ram[815]), .A(ram[831]), .S(n12679), .Y(n12508) );
  MUX2X1 U13022 ( .B(ram[783]), .A(ram[799]), .S(n12679), .Y(n12507) );
  MUX2X1 U13023 ( .B(n12506), .A(n12503), .S(n12585), .Y(n12510) );
  MUX2X1 U13024 ( .B(ram[751]), .A(ram[767]), .S(n12680), .Y(n12514) );
  MUX2X1 U13025 ( .B(ram[719]), .A(ram[735]), .S(n12680), .Y(n12513) );
  MUX2X1 U13026 ( .B(ram[687]), .A(ram[703]), .S(n12680), .Y(n12517) );
  MUX2X1 U13027 ( .B(ram[655]), .A(ram[671]), .S(n12680), .Y(n12516) );
  MUX2X1 U13028 ( .B(n12515), .A(n12512), .S(n12585), .Y(n12526) );
  MUX2X1 U13029 ( .B(ram[623]), .A(ram[639]), .S(n12680), .Y(n12520) );
  MUX2X1 U13030 ( .B(ram[591]), .A(ram[607]), .S(n12680), .Y(n12519) );
  MUX2X1 U13031 ( .B(ram[559]), .A(ram[575]), .S(n12680), .Y(n12523) );
  MUX2X1 U13032 ( .B(ram[527]), .A(ram[543]), .S(n12680), .Y(n12522) );
  MUX2X1 U13033 ( .B(n12521), .A(n12518), .S(n12585), .Y(n12525) );
  MUX2X1 U13034 ( .B(n12524), .A(n12509), .S(n12567), .Y(n12559) );
  MUX2X1 U13035 ( .B(ram[495]), .A(ram[511]), .S(n12680), .Y(n12529) );
  MUX2X1 U13036 ( .B(ram[463]), .A(ram[479]), .S(n12680), .Y(n12528) );
  MUX2X1 U13037 ( .B(ram[431]), .A(ram[447]), .S(n12680), .Y(n12532) );
  MUX2X1 U13038 ( .B(ram[399]), .A(ram[415]), .S(n12680), .Y(n12531) );
  MUX2X1 U13039 ( .B(n12530), .A(n12527), .S(n12585), .Y(n12541) );
  MUX2X1 U13040 ( .B(ram[367]), .A(ram[383]), .S(n12681), .Y(n12535) );
  MUX2X1 U13041 ( .B(ram[335]), .A(ram[351]), .S(n12681), .Y(n12534) );
  MUX2X1 U13042 ( .B(ram[303]), .A(ram[319]), .S(n12681), .Y(n12538) );
  MUX2X1 U13043 ( .B(ram[271]), .A(ram[287]), .S(n12681), .Y(n12537) );
  MUX2X1 U13044 ( .B(n12536), .A(n12533), .S(n12585), .Y(n12540) );
  MUX2X1 U13045 ( .B(ram[239]), .A(ram[255]), .S(n12681), .Y(n12544) );
  MUX2X1 U13046 ( .B(ram[207]), .A(ram[223]), .S(n12681), .Y(n12543) );
  MUX2X1 U13047 ( .B(ram[175]), .A(ram[191]), .S(n12681), .Y(n12547) );
  MUX2X1 U13048 ( .B(ram[143]), .A(ram[159]), .S(n12681), .Y(n12546) );
  MUX2X1 U13049 ( .B(n12545), .A(n12542), .S(n12585), .Y(n12556) );
  MUX2X1 U13050 ( .B(ram[111]), .A(ram[127]), .S(n12681), .Y(n12550) );
  MUX2X1 U13051 ( .B(ram[79]), .A(ram[95]), .S(n12681), .Y(n12549) );
  MUX2X1 U13052 ( .B(ram[47]), .A(ram[63]), .S(n12681), .Y(n12553) );
  MUX2X1 U13053 ( .B(ram[15]), .A(ram[31]), .S(n12681), .Y(n12552) );
  MUX2X1 U13054 ( .B(n12551), .A(n12548), .S(n12585), .Y(n12555) );
  MUX2X1 U13055 ( .B(n12554), .A(n12539), .S(n12567), .Y(n12558) );
  MUX2X1 U13056 ( .B(n12557), .A(n12494), .S(mem_access_addr[6]), .Y(n12560)
         );
  AND2X2 U13057 ( .A(n4384), .B(n4228), .Y(n324) );
  AND2X2 U13058 ( .A(n4384), .B(n4210), .Y(n306) );
  AND2X2 U13059 ( .A(n4384), .B(n4192), .Y(n288) );
  AND2X2 U13060 ( .A(n4384), .B(n4174), .Y(n270) );
  AND2X2 U13061 ( .A(n4315), .B(n4228), .Y(n252) );
  AND2X2 U13062 ( .A(n4315), .B(n4210), .Y(n234) );
  AND2X2 U13063 ( .A(n4315), .B(n4192), .Y(n216) );
  AND2X2 U13064 ( .A(n4315), .B(n4174), .Y(n198) );
  AND2X2 U13065 ( .A(n4246), .B(n4228), .Y(n180) );
  AND2X2 U13066 ( .A(n4246), .B(n4210), .Y(n162) );
  AND2X2 U13067 ( .A(n4246), .B(n4192), .Y(n144) );
  AND2X2 U13068 ( .A(n4246), .B(n4174), .Y(n126) );
  AND2X2 U13069 ( .A(n4228), .B(n4173), .Y(n108) );
  AND2X2 U13070 ( .A(n4210), .B(n4173), .Y(n90) );
  AND2X2 U13071 ( .A(n4192), .B(n4173), .Y(n72) );
  AND2X2 U13072 ( .A(n4173), .B(n4174), .Y(n54) );
  INVX2 U13073 ( .A(mem_write_data[15]), .Y(n13056) );
  INVX2 U13074 ( .A(mem_write_data[14]), .Y(n13057) );
  INVX2 U13075 ( .A(mem_write_data[13]), .Y(n13058) );
  INVX2 U13076 ( .A(mem_write_data[12]), .Y(n13059) );
  INVX2 U13077 ( .A(mem_write_data[11]), .Y(n13060) );
  INVX2 U13078 ( .A(mem_write_data[10]), .Y(n13061) );
  INVX2 U13079 ( .A(mem_write_data[9]), .Y(n13062) );
  INVX2 U13080 ( .A(mem_write_data[8]), .Y(n13063) );
  INVX2 U13081 ( .A(mem_write_data[7]), .Y(n13064) );
  INVX2 U13082 ( .A(mem_write_data[6]), .Y(n13065) );
  INVX2 U13083 ( .A(mem_write_data[5]), .Y(n13066) );
  INVX2 U13084 ( .A(mem_write_data[4]), .Y(n13067) );
  INVX2 U13085 ( .A(mem_write_data[3]), .Y(n13068) );
  INVX2 U13086 ( .A(mem_write_data[2]), .Y(n13069) );
  INVX2 U13087 ( .A(mem_write_data[1]), .Y(n13070) );
  INVX2 U13088 ( .A(mem_write_data[0]), .Y(n13071) );
endmodule


module MEM_stage ( clk, rst, pipeline_reg_in, pipeline_reg_out );
  input [38:0] pipeline_reg_in;
  output [37:0] pipeline_reg_out;
  input clk, rst;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, n1, n2, n3;
  wire   [15:0] mem_read_data;

  DFFPOSX1 pipeline_reg_out_reg_37_ ( .D(N40), .CLK(clk), .Q(
        pipeline_reg_out[37]) );
  DFFPOSX1 pipeline_reg_out_reg_36_ ( .D(N39), .CLK(clk), .Q(
        pipeline_reg_out[36]) );
  DFFPOSX1 pipeline_reg_out_reg_35_ ( .D(N38), .CLK(clk), .Q(
        pipeline_reg_out[35]) );
  DFFPOSX1 pipeline_reg_out_reg_34_ ( .D(N37), .CLK(clk), .Q(
        pipeline_reg_out[34]) );
  DFFPOSX1 pipeline_reg_out_reg_33_ ( .D(N36), .CLK(clk), .Q(
        pipeline_reg_out[33]) );
  DFFPOSX1 pipeline_reg_out_reg_32_ ( .D(N35), .CLK(clk), .Q(
        pipeline_reg_out[32]) );
  DFFPOSX1 pipeline_reg_out_reg_31_ ( .D(N34), .CLK(clk), .Q(
        pipeline_reg_out[31]) );
  DFFPOSX1 pipeline_reg_out_reg_30_ ( .D(N33), .CLK(clk), .Q(
        pipeline_reg_out[30]) );
  DFFPOSX1 pipeline_reg_out_reg_29_ ( .D(N32), .CLK(clk), .Q(
        pipeline_reg_out[29]) );
  DFFPOSX1 pipeline_reg_out_reg_28_ ( .D(N31), .CLK(clk), .Q(
        pipeline_reg_out[28]) );
  DFFPOSX1 pipeline_reg_out_reg_27_ ( .D(N30), .CLK(clk), .Q(
        pipeline_reg_out[27]) );
  DFFPOSX1 pipeline_reg_out_reg_26_ ( .D(N29), .CLK(clk), .Q(
        pipeline_reg_out[26]) );
  DFFPOSX1 pipeline_reg_out_reg_25_ ( .D(N28), .CLK(clk), .Q(
        pipeline_reg_out[25]) );
  DFFPOSX1 pipeline_reg_out_reg_24_ ( .D(N27), .CLK(clk), .Q(
        pipeline_reg_out[24]) );
  DFFPOSX1 pipeline_reg_out_reg_23_ ( .D(N26), .CLK(clk), .Q(
        pipeline_reg_out[23]) );
  DFFPOSX1 pipeline_reg_out_reg_22_ ( .D(N25), .CLK(clk), .Q(
        pipeline_reg_out[22]) );
  DFFPOSX1 pipeline_reg_out_reg_21_ ( .D(N24), .CLK(clk), .Q(
        pipeline_reg_out[21]) );
  DFFPOSX1 pipeline_reg_out_reg_20_ ( .D(N23), .CLK(clk), .Q(
        pipeline_reg_out[20]) );
  DFFPOSX1 pipeline_reg_out_reg_19_ ( .D(N22), .CLK(clk), .Q(
        pipeline_reg_out[19]) );
  DFFPOSX1 pipeline_reg_out_reg_18_ ( .D(N21), .CLK(clk), .Q(
        pipeline_reg_out[18]) );
  DFFPOSX1 pipeline_reg_out_reg_17_ ( .D(N20), .CLK(clk), .Q(
        pipeline_reg_out[17]) );
  DFFPOSX1 pipeline_reg_out_reg_16_ ( .D(N19), .CLK(clk), .Q(
        pipeline_reg_out[16]) );
  DFFPOSX1 pipeline_reg_out_reg_15_ ( .D(N18), .CLK(clk), .Q(
        pipeline_reg_out[15]) );
  DFFPOSX1 pipeline_reg_out_reg_14_ ( .D(N17), .CLK(clk), .Q(
        pipeline_reg_out[14]) );
  DFFPOSX1 pipeline_reg_out_reg_13_ ( .D(N16), .CLK(clk), .Q(
        pipeline_reg_out[13]) );
  DFFPOSX1 pipeline_reg_out_reg_12_ ( .D(N15), .CLK(clk), .Q(
        pipeline_reg_out[12]) );
  DFFPOSX1 pipeline_reg_out_reg_11_ ( .D(N14), .CLK(clk), .Q(
        pipeline_reg_out[11]) );
  DFFPOSX1 pipeline_reg_out_reg_10_ ( .D(N13), .CLK(clk), .Q(
        pipeline_reg_out[10]) );
  DFFPOSX1 pipeline_reg_out_reg_9_ ( .D(N12), .CLK(clk), .Q(
        pipeline_reg_out[9]) );
  DFFPOSX1 pipeline_reg_out_reg_8_ ( .D(N11), .CLK(clk), .Q(
        pipeline_reg_out[8]) );
  DFFPOSX1 pipeline_reg_out_reg_7_ ( .D(N10), .CLK(clk), .Q(
        pipeline_reg_out[7]) );
  DFFPOSX1 pipeline_reg_out_reg_6_ ( .D(N9), .CLK(clk), .Q(pipeline_reg_out[6]) );
  DFFPOSX1 pipeline_reg_out_reg_5_ ( .D(N8), .CLK(clk), .Q(pipeline_reg_out[5]) );
  DFFPOSX1 pipeline_reg_out_reg_4_ ( .D(N7), .CLK(clk), .Q(pipeline_reg_out[4]) );
  DFFPOSX1 pipeline_reg_out_reg_3_ ( .D(N6), .CLK(clk), .Q(pipeline_reg_out[3]) );
  DFFPOSX1 pipeline_reg_out_reg_2_ ( .D(N5), .CLK(clk), .Q(pipeline_reg_out[2]) );
  DFFPOSX1 pipeline_reg_out_reg_1_ ( .D(N4), .CLK(clk), .Q(pipeline_reg_out[1]) );
  DFFPOSX1 pipeline_reg_out_reg_0_ ( .D(N3), .CLK(clk), .Q(pipeline_reg_out[0]) );
  AND2X1 U4 ( .A(mem_read_data[1]), .B(n3), .Y(N9) );
  AND2X1 U5 ( .A(mem_read_data[0]), .B(n3), .Y(N8) );
  AND2X1 U6 ( .A(pipeline_reg_in[4]), .B(n3), .Y(N7) );
  AND2X1 U7 ( .A(pipeline_reg_in[3]), .B(n3), .Y(N6) );
  AND2X1 U8 ( .A(pipeline_reg_in[2]), .B(n3), .Y(N5) );
  AND2X1 U9 ( .A(pipeline_reg_in[38]), .B(n3), .Y(N40) );
  AND2X1 U10 ( .A(pipeline_reg_in[1]), .B(n3), .Y(N4) );
  AND2X1 U11 ( .A(pipeline_reg_in[37]), .B(n3), .Y(N39) );
  AND2X1 U12 ( .A(pipeline_reg_in[36]), .B(n3), .Y(N38) );
  AND2X1 U13 ( .A(pipeline_reg_in[35]), .B(n3), .Y(N37) );
  AND2X1 U14 ( .A(pipeline_reg_in[34]), .B(n3), .Y(N36) );
  AND2X1 U15 ( .A(pipeline_reg_in[33]), .B(n3), .Y(N35) );
  AND2X1 U16 ( .A(pipeline_reg_in[32]), .B(n3), .Y(N34) );
  AND2X1 U17 ( .A(pipeline_reg_in[31]), .B(n3), .Y(N33) );
  AND2X1 U18 ( .A(pipeline_reg_in[30]), .B(n3), .Y(N32) );
  AND2X1 U19 ( .A(pipeline_reg_in[29]), .B(n3), .Y(N31) );
  AND2X1 U20 ( .A(pipeline_reg_in[28]), .B(n3), .Y(N30) );
  AND2X1 U21 ( .A(pipeline_reg_in[0]), .B(n3), .Y(N3) );
  AND2X1 U22 ( .A(pipeline_reg_in[27]), .B(n3), .Y(N29) );
  AND2X1 U23 ( .A(pipeline_reg_in[26]), .B(n3), .Y(N28) );
  AND2X1 U24 ( .A(n1), .B(n3), .Y(N27) );
  AND2X1 U25 ( .A(pipeline_reg_in[24]), .B(n3), .Y(N26) );
  AND2X1 U26 ( .A(pipeline_reg_in[23]), .B(n3), .Y(N25) );
  AND2X1 U27 ( .A(pipeline_reg_in[22]), .B(n3), .Y(N24) );
  AND2X1 U28 ( .A(mem_read_data[15]), .B(n3), .Y(N23) );
  AND2X1 U29 ( .A(mem_read_data[14]), .B(n3), .Y(N22) );
  AND2X1 U30 ( .A(mem_read_data[13]), .B(n3), .Y(N21) );
  AND2X1 U31 ( .A(mem_read_data[12]), .B(n3), .Y(N20) );
  AND2X1 U32 ( .A(mem_read_data[11]), .B(n3), .Y(N19) );
  AND2X1 U33 ( .A(mem_read_data[10]), .B(n3), .Y(N18) );
  AND2X1 U34 ( .A(mem_read_data[9]), .B(n3), .Y(N17) );
  AND2X1 U35 ( .A(mem_read_data[8]), .B(n3), .Y(N16) );
  AND2X1 U36 ( .A(mem_read_data[7]), .B(n3), .Y(N15) );
  AND2X1 U37 ( .A(mem_read_data[6]), .B(n3), .Y(N14) );
  AND2X1 U38 ( .A(mem_read_data[5]), .B(n3), .Y(N13) );
  AND2X1 U39 ( .A(mem_read_data[4]), .B(n3), .Y(N12) );
  AND2X1 U40 ( .A(mem_read_data[3]), .B(n3), .Y(N11) );
  AND2X1 U41 ( .A(mem_read_data[2]), .B(n3), .Y(N10) );
  data_mem dmem ( .clk(clk), .mem_access_addr({pipeline_reg_in[37:26], n1, 
        pipeline_reg_in[24:22]}), .mem_write_data(pipeline_reg_in[20:5]), 
        .mem_write_en(pipeline_reg_in[21]), .mem_read_data(mem_read_data) );
  INVX2 U3 ( .A(n2), .Y(n1) );
  INVX2 U42 ( .A(pipeline_reg_in[25]), .Y(n2) );
  INVX2 U43 ( .A(rst), .Y(n3) );
endmodule


module WB_stage ( clk, rst, pipeline_reg_in, reg_write_en, reg_write_dest, 
        reg_write_data, instruction_fetch_en );
  input [37:0] pipeline_reg_in;
  output [2:0] reg_write_dest;
  output [15:0] reg_write_data;
  input clk, rst;
  output reg_write_en, instruction_fetch_en;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n1, n20, n22, n24, n26, n27;

  DFFSR instruction_fetch_en_reg ( .D(pipeline_reg_in[37]), .CLK(clk), .R(1'b1), .S(n27), .Q(instruction_fetch_en) );
  INVX2 U5 ( .A(n4), .Y(reg_write_data[9]) );
  INVX2 U6 ( .A(n5), .Y(reg_write_data[8]) );
  INVX2 U7 ( .A(n6), .Y(reg_write_data[7]) );
  INVX2 U8 ( .A(n7), .Y(reg_write_data[6]) );
  INVX2 U9 ( .A(n8), .Y(reg_write_data[5]) );
  INVX2 U10 ( .A(n9), .Y(reg_write_data[4]) );
  INVX2 U11 ( .A(n10), .Y(reg_write_data[3]) );
  INVX2 U12 ( .A(n11), .Y(reg_write_data[2]) );
  INVX2 U13 ( .A(n12), .Y(reg_write_data[1]) );
  INVX2 U14 ( .A(n13), .Y(reg_write_data[15]) );
  INVX2 U15 ( .A(n14), .Y(reg_write_data[14]) );
  INVX2 U16 ( .A(n15), .Y(reg_write_data[13]) );
  INVX2 U17 ( .A(n16), .Y(reg_write_data[12]) );
  INVX2 U18 ( .A(n17), .Y(reg_write_data[11]) );
  INVX2 U19 ( .A(n18), .Y(reg_write_data[10]) );
  INVX2 U20 ( .A(n19), .Y(reg_write_data[0]) );
  AOI22X1 U22 ( .A(pipeline_reg_in[0]), .B(pipeline_reg_in[14]), .C(
        pipeline_reg_in[30]), .D(n26), .Y(n4) );
  AOI22X1 U23 ( .A(pipeline_reg_in[13]), .B(pipeline_reg_in[0]), .C(
        pipeline_reg_in[29]), .D(n26), .Y(n5) );
  AOI22X1 U24 ( .A(pipeline_reg_in[12]), .B(pipeline_reg_in[0]), .C(
        pipeline_reg_in[28]), .D(n26), .Y(n6) );
  AOI22X1 U25 ( .A(pipeline_reg_in[11]), .B(pipeline_reg_in[0]), .C(
        pipeline_reg_in[27]), .D(n26), .Y(n7) );
  AOI22X1 U26 ( .A(pipeline_reg_in[10]), .B(pipeline_reg_in[0]), .C(
        pipeline_reg_in[26]), .D(n26), .Y(n8) );
  AOI22X1 U27 ( .A(pipeline_reg_in[25]), .B(n26), .C(pipeline_reg_in[9]), .D(
        pipeline_reg_in[0]), .Y(n9) );
  AOI22X1 U28 ( .A(pipeline_reg_in[24]), .B(n26), .C(pipeline_reg_in[8]), .D(
        pipeline_reg_in[0]), .Y(n10) );
  AOI22X1 U29 ( .A(pipeline_reg_in[23]), .B(n26), .C(pipeline_reg_in[7]), .D(
        pipeline_reg_in[0]), .Y(n11) );
  AOI22X1 U30 ( .A(pipeline_reg_in[22]), .B(n26), .C(pipeline_reg_in[6]), .D(
        pipeline_reg_in[0]), .Y(n12) );
  AOI22X1 U31 ( .A(pipeline_reg_in[20]), .B(pipeline_reg_in[0]), .C(
        pipeline_reg_in[36]), .D(n26), .Y(n13) );
  AOI22X1 U32 ( .A(pipeline_reg_in[19]), .B(pipeline_reg_in[0]), .C(
        pipeline_reg_in[35]), .D(n26), .Y(n14) );
  AOI22X1 U33 ( .A(pipeline_reg_in[18]), .B(pipeline_reg_in[0]), .C(
        pipeline_reg_in[34]), .D(n26), .Y(n15) );
  AOI22X1 U34 ( .A(pipeline_reg_in[17]), .B(pipeline_reg_in[0]), .C(
        pipeline_reg_in[33]), .D(n26), .Y(n16) );
  AOI22X1 U35 ( .A(pipeline_reg_in[16]), .B(pipeline_reg_in[0]), .C(
        pipeline_reg_in[32]), .D(n26), .Y(n17) );
  AOI22X1 U36 ( .A(pipeline_reg_in[15]), .B(pipeline_reg_in[0]), .C(
        pipeline_reg_in[31]), .D(n26), .Y(n18) );
  AOI22X1 U37 ( .A(pipeline_reg_in[21]), .B(n26), .C(pipeline_reg_in[5]), .D(
        pipeline_reg_in[0]), .Y(n19) );
  INVX2 U3 ( .A(pipeline_reg_in[0]), .Y(n26) );
  INVX2 U21 ( .A(n24), .Y(reg_write_en) );
  INVX2 U38 ( .A(pipeline_reg_in[4]), .Y(n24) );
  INVX2 U39 ( .A(n22), .Y(reg_write_dest[2]) );
  INVX2 U40 ( .A(pipeline_reg_in[3]), .Y(n22) );
  INVX2 U41 ( .A(n20), .Y(reg_write_dest[1]) );
  INVX2 U42 ( .A(pipeline_reg_in[2]), .Y(n20) );
  INVX2 U43 ( .A(n1), .Y(reg_write_dest[0]) );
  INVX2 U44 ( .A(pipeline_reg_in[1]), .Y(n1) );
  INVX2 U45 ( .A(rst), .Y(n27) );
endmodule


module register_file ( clk, rst, reg_write_en, reg_write_dest, reg_write_data, 
        reg_read_addr_1, reg_read_data_1, reg_read_addr_2, reg_read_data_2 );
  input [2:0] reg_write_dest;
  input [15:0] reg_write_data;
  input [2:0] reg_read_addr_1;
  output [15:0] reg_read_data_1;
  input [2:0] reg_read_addr_2;
  output [15:0] reg_read_data_2;
  input clk, rst, reg_write_en;
  wire   N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42,
         N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N59, N60, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n128, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671;
  wire   [127:0] reg_array;

  DFFSR reg_array_reg_7__15_ ( .D(n418), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[127]) );
  DFFSR reg_array_reg_7__14_ ( .D(n417), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[126]) );
  DFFSR reg_array_reg_7__13_ ( .D(n416), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[125]) );
  DFFSR reg_array_reg_7__12_ ( .D(n415), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[124]) );
  DFFSR reg_array_reg_7__11_ ( .D(n414), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[123]) );
  DFFSR reg_array_reg_7__10_ ( .D(n413), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[122]) );
  DFFSR reg_array_reg_7__9_ ( .D(n412), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[121]) );
  DFFSR reg_array_reg_7__8_ ( .D(n411), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[120]) );
  DFFSR reg_array_reg_7__7_ ( .D(n410), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[119]) );
  DFFSR reg_array_reg_7__6_ ( .D(n409), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[118]) );
  DFFSR reg_array_reg_7__5_ ( .D(n408), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[117]) );
  DFFSR reg_array_reg_7__4_ ( .D(n407), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[116]) );
  DFFSR reg_array_reg_7__3_ ( .D(n406), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[115]) );
  DFFSR reg_array_reg_7__2_ ( .D(n405), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[114]) );
  DFFSR reg_array_reg_7__1_ ( .D(n404), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[113]) );
  DFFSR reg_array_reg_7__0_ ( .D(n403), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[112]) );
  DFFSR reg_array_reg_6__15_ ( .D(n402), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[111]) );
  DFFSR reg_array_reg_6__14_ ( .D(n401), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[110]) );
  DFFSR reg_array_reg_6__13_ ( .D(n400), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[109]) );
  DFFSR reg_array_reg_6__12_ ( .D(n399), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[108]) );
  DFFSR reg_array_reg_6__11_ ( .D(n398), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[107]) );
  DFFSR reg_array_reg_6__10_ ( .D(n397), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[106]) );
  DFFSR reg_array_reg_6__9_ ( .D(n396), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[105]) );
  DFFSR reg_array_reg_6__8_ ( .D(n395), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[104]) );
  DFFSR reg_array_reg_6__7_ ( .D(n394), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[103]) );
  DFFSR reg_array_reg_6__6_ ( .D(n393), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[102]) );
  DFFSR reg_array_reg_6__5_ ( .D(n392), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[101]) );
  DFFSR reg_array_reg_6__4_ ( .D(n391), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[100]) );
  DFFSR reg_array_reg_6__3_ ( .D(n390), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[99]) );
  DFFSR reg_array_reg_6__2_ ( .D(n389), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[98]) );
  DFFSR reg_array_reg_6__1_ ( .D(n388), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[97]) );
  DFFSR reg_array_reg_6__0_ ( .D(n387), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[96]) );
  DFFSR reg_array_reg_5__15_ ( .D(n386), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[95]) );
  DFFSR reg_array_reg_5__14_ ( .D(n385), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[94]) );
  DFFSR reg_array_reg_5__13_ ( .D(n384), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[93]) );
  DFFSR reg_array_reg_5__12_ ( .D(n383), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[92]) );
  DFFSR reg_array_reg_5__11_ ( .D(n382), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[91]) );
  DFFSR reg_array_reg_5__10_ ( .D(n381), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[90]) );
  DFFSR reg_array_reg_5__9_ ( .D(n380), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[89]) );
  DFFSR reg_array_reg_5__8_ ( .D(n379), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[88]) );
  DFFSR reg_array_reg_5__7_ ( .D(n378), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[87]) );
  DFFSR reg_array_reg_5__6_ ( .D(n377), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[86]) );
  DFFSR reg_array_reg_5__5_ ( .D(n376), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[85]) );
  DFFSR reg_array_reg_5__4_ ( .D(n375), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[84]) );
  DFFSR reg_array_reg_5__3_ ( .D(n374), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[83]) );
  DFFSR reg_array_reg_5__2_ ( .D(n373), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[82]) );
  DFFSR reg_array_reg_5__1_ ( .D(n372), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[81]) );
  DFFSR reg_array_reg_5__0_ ( .D(n371), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[80]) );
  DFFSR reg_array_reg_4__15_ ( .D(n370), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[79]) );
  DFFSR reg_array_reg_4__14_ ( .D(n369), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[78]) );
  DFFSR reg_array_reg_4__13_ ( .D(n368), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[77]) );
  DFFSR reg_array_reg_4__12_ ( .D(n367), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[76]) );
  DFFSR reg_array_reg_4__11_ ( .D(n366), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[75]) );
  DFFSR reg_array_reg_4__10_ ( .D(n365), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[74]) );
  DFFSR reg_array_reg_4__9_ ( .D(n364), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[73]) );
  DFFSR reg_array_reg_4__8_ ( .D(n363), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[72]) );
  DFFSR reg_array_reg_4__7_ ( .D(n362), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[71]) );
  DFFSR reg_array_reg_4__6_ ( .D(n361), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[70]) );
  DFFSR reg_array_reg_4__5_ ( .D(n360), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[69]) );
  DFFSR reg_array_reg_4__4_ ( .D(n359), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[68]) );
  DFFSR reg_array_reg_4__3_ ( .D(n358), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[67]) );
  DFFSR reg_array_reg_4__2_ ( .D(n357), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[66]) );
  DFFSR reg_array_reg_4__1_ ( .D(n356), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[65]) );
  DFFSR reg_array_reg_4__0_ ( .D(n355), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[64]) );
  DFFSR reg_array_reg_3__15_ ( .D(n354), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[63]) );
  DFFSR reg_array_reg_3__14_ ( .D(n353), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[62]) );
  DFFSR reg_array_reg_3__13_ ( .D(n352), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[61]) );
  DFFSR reg_array_reg_3__12_ ( .D(n351), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[60]) );
  DFFSR reg_array_reg_3__11_ ( .D(n350), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[59]) );
  DFFSR reg_array_reg_3__10_ ( .D(n349), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[58]) );
  DFFSR reg_array_reg_3__9_ ( .D(n348), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[57]) );
  DFFSR reg_array_reg_3__8_ ( .D(n347), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[56]) );
  DFFSR reg_array_reg_3__7_ ( .D(n346), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[55]) );
  DFFSR reg_array_reg_3__6_ ( .D(n345), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[54]) );
  DFFSR reg_array_reg_3__5_ ( .D(n344), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[53]) );
  DFFSR reg_array_reg_3__4_ ( .D(n343), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[52]) );
  DFFSR reg_array_reg_3__3_ ( .D(n342), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[51]) );
  DFFSR reg_array_reg_3__2_ ( .D(n341), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[50]) );
  DFFSR reg_array_reg_3__1_ ( .D(n340), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[49]) );
  DFFSR reg_array_reg_3__0_ ( .D(n339), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[48]) );
  DFFSR reg_array_reg_2__15_ ( .D(n338), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[47]) );
  DFFSR reg_array_reg_2__14_ ( .D(n337), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[46]) );
  DFFSR reg_array_reg_2__13_ ( .D(n336), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[45]) );
  DFFSR reg_array_reg_2__12_ ( .D(n335), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[44]) );
  DFFSR reg_array_reg_2__11_ ( .D(n334), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[43]) );
  DFFSR reg_array_reg_2__10_ ( .D(n333), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[42]) );
  DFFSR reg_array_reg_2__9_ ( .D(n332), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[41]) );
  DFFSR reg_array_reg_2__8_ ( .D(n331), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[40]) );
  DFFSR reg_array_reg_2__7_ ( .D(n330), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[39]) );
  DFFSR reg_array_reg_2__6_ ( .D(n329), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[38]) );
  DFFSR reg_array_reg_2__5_ ( .D(n328), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[37]) );
  DFFSR reg_array_reg_2__4_ ( .D(n327), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[36]) );
  DFFSR reg_array_reg_2__3_ ( .D(n326), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[35]) );
  DFFSR reg_array_reg_2__2_ ( .D(n325), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[34]) );
  DFFSR reg_array_reg_2__1_ ( .D(n324), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[33]) );
  DFFSR reg_array_reg_2__0_ ( .D(n323), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[32]) );
  DFFSR reg_array_reg_1__15_ ( .D(n322), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[31]) );
  DFFSR reg_array_reg_1__14_ ( .D(n321), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[30]) );
  DFFSR reg_array_reg_1__13_ ( .D(n320), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[29]) );
  DFFSR reg_array_reg_1__12_ ( .D(n319), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[28]) );
  DFFSR reg_array_reg_1__11_ ( .D(n318), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[27]) );
  DFFSR reg_array_reg_1__10_ ( .D(n317), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[26]) );
  DFFSR reg_array_reg_1__9_ ( .D(n316), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[25]) );
  DFFSR reg_array_reg_1__8_ ( .D(n315), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[24]) );
  DFFSR reg_array_reg_1__7_ ( .D(n314), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[23]) );
  DFFSR reg_array_reg_1__6_ ( .D(n313), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[22]) );
  DFFSR reg_array_reg_1__5_ ( .D(n312), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[21]) );
  DFFSR reg_array_reg_1__4_ ( .D(n311), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[20]) );
  DFFSR reg_array_reg_1__3_ ( .D(n310), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[19]) );
  DFFSR reg_array_reg_1__2_ ( .D(n309), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[18]) );
  DFFSR reg_array_reg_1__1_ ( .D(n308), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[17]) );
  DFFSR reg_array_reg_1__0_ ( .D(n307), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[16]) );
  DFFSR reg_array_reg_0__15_ ( .D(n306), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[15]) );
  DFFSR reg_array_reg_0__14_ ( .D(n305), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[14]) );
  DFFSR reg_array_reg_0__13_ ( .D(n304), .CLK(clk), .R(n633), .S(1'b1), .Q(
        reg_array[13]) );
  DFFSR reg_array_reg_0__12_ ( .D(n303), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[12]) );
  DFFSR reg_array_reg_0__11_ ( .D(n302), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[11]) );
  DFFSR reg_array_reg_0__10_ ( .D(n301), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[10]) );
  DFFSR reg_array_reg_0__9_ ( .D(n300), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[9]) );
  DFFSR reg_array_reg_0__8_ ( .D(n299), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[8]) );
  DFFSR reg_array_reg_0__7_ ( .D(n298), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[7]) );
  DFFSR reg_array_reg_0__6_ ( .D(n297), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[6]) );
  DFFSR reg_array_reg_0__5_ ( .D(n296), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[5]) );
  DFFSR reg_array_reg_0__4_ ( .D(n295), .CLK(clk), .R(n632), .S(1'b1), .Q(
        reg_array[4]) );
  DFFSR reg_array_reg_0__3_ ( .D(n294), .CLK(clk), .R(n630), .S(1'b1), .Q(
        reg_array[3]) );
  DFFSR reg_array_reg_0__2_ ( .D(n293), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[2]) );
  DFFSR reg_array_reg_0__1_ ( .D(n292), .CLK(clk), .R(n671), .S(1'b1), .Q(
        reg_array[1]) );
  DFFSR reg_array_reg_0__0_ ( .D(n291), .CLK(clk), .R(n631), .S(1'b1), .Q(
        reg_array[0]) );
  AND2X1 U152 ( .A(N51), .B(n669), .Y(reg_read_data_2[9]) );
  AND2X1 U153 ( .A(N52), .B(n669), .Y(reg_read_data_2[8]) );
  AND2X1 U154 ( .A(N53), .B(n669), .Y(reg_read_data_2[7]) );
  AND2X1 U155 ( .A(N54), .B(n669), .Y(reg_read_data_2[6]) );
  AND2X1 U156 ( .A(N55), .B(n669), .Y(reg_read_data_2[5]) );
  AND2X1 U157 ( .A(N56), .B(n669), .Y(reg_read_data_2[4]) );
  AND2X1 U158 ( .A(N57), .B(n669), .Y(reg_read_data_2[3]) );
  AND2X1 U159 ( .A(N58), .B(n669), .Y(reg_read_data_2[2]) );
  AND2X1 U160 ( .A(N59), .B(n669), .Y(reg_read_data_2[1]) );
  AND2X1 U161 ( .A(N45), .B(n669), .Y(reg_read_data_2[15]) );
  AND2X1 U162 ( .A(N46), .B(n669), .Y(reg_read_data_2[14]) );
  AND2X1 U163 ( .A(N47), .B(n669), .Y(reg_read_data_2[13]) );
  AND2X1 U164 ( .A(N48), .B(n669), .Y(reg_read_data_2[12]) );
  AND2X1 U165 ( .A(N49), .B(n669), .Y(reg_read_data_2[11]) );
  AND2X1 U166 ( .A(N50), .B(n669), .Y(reg_read_data_2[10]) );
  AND2X1 U167 ( .A(N60), .B(n669), .Y(reg_read_data_2[0]) );
  NOR3X1 U168 ( .A(reg_read_addr_2[1]), .B(reg_read_addr_2[2]), .C(
        reg_read_addr_2[0]), .Y(n151) );
  AND2X1 U169 ( .A(N35), .B(n670), .Y(reg_read_data_1[9]) );
  AND2X1 U170 ( .A(N36), .B(n670), .Y(reg_read_data_1[8]) );
  AND2X1 U171 ( .A(N37), .B(n670), .Y(reg_read_data_1[7]) );
  AND2X1 U172 ( .A(N38), .B(n670), .Y(reg_read_data_1[6]) );
  AND2X1 U173 ( .A(N39), .B(n670), .Y(reg_read_data_1[5]) );
  AND2X1 U174 ( .A(N40), .B(n670), .Y(reg_read_data_1[4]) );
  AND2X1 U175 ( .A(N41), .B(n670), .Y(reg_read_data_1[3]) );
  AND2X1 U176 ( .A(N42), .B(n670), .Y(reg_read_data_1[2]) );
  AND2X1 U177 ( .A(N43), .B(n670), .Y(reg_read_data_1[1]) );
  AND2X1 U178 ( .A(N29), .B(n670), .Y(reg_read_data_1[15]) );
  AND2X1 U179 ( .A(N30), .B(n670), .Y(reg_read_data_1[14]) );
  AND2X1 U180 ( .A(N31), .B(n670), .Y(reg_read_data_1[13]) );
  AND2X1 U181 ( .A(N32), .B(n670), .Y(reg_read_data_1[12]) );
  AND2X1 U182 ( .A(N33), .B(n670), .Y(reg_read_data_1[11]) );
  AND2X1 U183 ( .A(N34), .B(n670), .Y(reg_read_data_1[10]) );
  AND2X1 U184 ( .A(N44), .B(n670), .Y(reg_read_data_1[0]) );
  NOR3X1 U185 ( .A(n128), .B(reg_read_addr_1[2]), .C(reg_read_addr_1[0]), .Y(
        n152) );
  OAI21X1 U186 ( .A(n648), .B(n665), .C(n154), .Y(n291) );
  NAND2X1 U187 ( .A(reg_array[0]), .B(n648), .Y(n154) );
  OAI21X1 U188 ( .A(n648), .B(n664), .C(n155), .Y(n292) );
  NAND2X1 U189 ( .A(reg_array[1]), .B(n648), .Y(n155) );
  OAI21X1 U190 ( .A(n648), .B(n663), .C(n156), .Y(n293) );
  NAND2X1 U191 ( .A(reg_array[2]), .B(n153), .Y(n156) );
  OAI21X1 U192 ( .A(n648), .B(n662), .C(n157), .Y(n294) );
  NAND2X1 U193 ( .A(reg_array[3]), .B(n153), .Y(n157) );
  OAI21X1 U194 ( .A(n648), .B(n661), .C(n158), .Y(n295) );
  NAND2X1 U195 ( .A(reg_array[4]), .B(n153), .Y(n158) );
  OAI21X1 U196 ( .A(n648), .B(n660), .C(n159), .Y(n296) );
  NAND2X1 U197 ( .A(reg_array[5]), .B(n153), .Y(n159) );
  OAI21X1 U198 ( .A(n648), .B(n659), .C(n160), .Y(n297) );
  NAND2X1 U199 ( .A(reg_array[6]), .B(n153), .Y(n160) );
  OAI21X1 U200 ( .A(n648), .B(n658), .C(n161), .Y(n298) );
  NAND2X1 U201 ( .A(reg_array[7]), .B(n153), .Y(n161) );
  OAI21X1 U202 ( .A(n648), .B(n657), .C(n162), .Y(n299) );
  NAND2X1 U203 ( .A(reg_array[8]), .B(n153), .Y(n162) );
  OAI21X1 U204 ( .A(n648), .B(n656), .C(n163), .Y(n300) );
  NAND2X1 U205 ( .A(reg_array[9]), .B(n153), .Y(n163) );
  OAI21X1 U206 ( .A(n648), .B(n655), .C(n164), .Y(n301) );
  NAND2X1 U207 ( .A(reg_array[10]), .B(n153), .Y(n164) );
  OAI21X1 U208 ( .A(n648), .B(n654), .C(n165), .Y(n302) );
  NAND2X1 U209 ( .A(reg_array[11]), .B(n153), .Y(n165) );
  OAI21X1 U210 ( .A(n153), .B(n653), .C(n166), .Y(n303) );
  NAND2X1 U211 ( .A(reg_array[12]), .B(n153), .Y(n166) );
  OAI21X1 U212 ( .A(n153), .B(n652), .C(n167), .Y(n304) );
  NAND2X1 U213 ( .A(reg_array[13]), .B(n153), .Y(n167) );
  OAI21X1 U214 ( .A(n153), .B(n651), .C(n168), .Y(n305) );
  NAND2X1 U215 ( .A(reg_array[14]), .B(n648), .Y(n168) );
  OAI21X1 U216 ( .A(n153), .B(n650), .C(n169), .Y(n306) );
  NAND2X1 U217 ( .A(reg_array[15]), .B(n648), .Y(n169) );
  NAND3X1 U218 ( .A(n668), .B(n667), .C(n170), .Y(n153) );
  OAI21X1 U219 ( .A(n665), .B(n646), .C(n172), .Y(n307) );
  NAND2X1 U220 ( .A(reg_array[16]), .B(n646), .Y(n172) );
  OAI21X1 U221 ( .A(n664), .B(n646), .C(n173), .Y(n308) );
  NAND2X1 U222 ( .A(reg_array[17]), .B(n646), .Y(n173) );
  OAI21X1 U223 ( .A(n663), .B(n646), .C(n174), .Y(n309) );
  NAND2X1 U224 ( .A(reg_array[18]), .B(n171), .Y(n174) );
  OAI21X1 U225 ( .A(n662), .B(n646), .C(n175), .Y(n310) );
  NAND2X1 U226 ( .A(reg_array[19]), .B(n171), .Y(n175) );
  OAI21X1 U227 ( .A(n661), .B(n646), .C(n176), .Y(n311) );
  NAND2X1 U228 ( .A(reg_array[20]), .B(n171), .Y(n176) );
  OAI21X1 U229 ( .A(n660), .B(n646), .C(n177), .Y(n312) );
  NAND2X1 U230 ( .A(reg_array[21]), .B(n171), .Y(n177) );
  OAI21X1 U231 ( .A(n659), .B(n646), .C(n178), .Y(n313) );
  NAND2X1 U232 ( .A(reg_array[22]), .B(n171), .Y(n178) );
  OAI21X1 U233 ( .A(n658), .B(n646), .C(n179), .Y(n314) );
  NAND2X1 U234 ( .A(reg_array[23]), .B(n171), .Y(n179) );
  OAI21X1 U235 ( .A(n657), .B(n646), .C(n180), .Y(n315) );
  NAND2X1 U236 ( .A(reg_array[24]), .B(n171), .Y(n180) );
  OAI21X1 U237 ( .A(n656), .B(n646), .C(n181), .Y(n316) );
  NAND2X1 U238 ( .A(reg_array[25]), .B(n171), .Y(n181) );
  OAI21X1 U239 ( .A(n655), .B(n646), .C(n182), .Y(n317) );
  NAND2X1 U240 ( .A(reg_array[26]), .B(n171), .Y(n182) );
  OAI21X1 U241 ( .A(n654), .B(n646), .C(n183), .Y(n318) );
  NAND2X1 U242 ( .A(reg_array[27]), .B(n171), .Y(n183) );
  OAI21X1 U243 ( .A(n653), .B(n171), .C(n184), .Y(n319) );
  NAND2X1 U244 ( .A(reg_array[28]), .B(n171), .Y(n184) );
  OAI21X1 U245 ( .A(n652), .B(n171), .C(n185), .Y(n320) );
  NAND2X1 U246 ( .A(reg_array[29]), .B(n171), .Y(n185) );
  OAI21X1 U247 ( .A(n651), .B(n171), .C(n186), .Y(n321) );
  NAND2X1 U248 ( .A(reg_array[30]), .B(n646), .Y(n186) );
  OAI21X1 U249 ( .A(n650), .B(n171), .C(n187), .Y(n322) );
  NAND2X1 U250 ( .A(reg_array[31]), .B(n646), .Y(n187) );
  NAND3X1 U251 ( .A(n170), .B(n667), .C(reg_write_dest[0]), .Y(n171) );
  OAI21X1 U252 ( .A(n665), .B(n644), .C(n189), .Y(n323) );
  NAND2X1 U253 ( .A(reg_array[32]), .B(n644), .Y(n189) );
  OAI21X1 U254 ( .A(n664), .B(n644), .C(n190), .Y(n324) );
  NAND2X1 U255 ( .A(reg_array[33]), .B(n644), .Y(n190) );
  OAI21X1 U256 ( .A(n663), .B(n644), .C(n191), .Y(n325) );
  NAND2X1 U257 ( .A(reg_array[34]), .B(n188), .Y(n191) );
  OAI21X1 U258 ( .A(n662), .B(n644), .C(n192), .Y(n326) );
  NAND2X1 U259 ( .A(reg_array[35]), .B(n188), .Y(n192) );
  OAI21X1 U260 ( .A(n661), .B(n644), .C(n193), .Y(n327) );
  NAND2X1 U261 ( .A(reg_array[36]), .B(n188), .Y(n193) );
  OAI21X1 U262 ( .A(n660), .B(n644), .C(n194), .Y(n328) );
  NAND2X1 U263 ( .A(reg_array[37]), .B(n188), .Y(n194) );
  OAI21X1 U264 ( .A(n659), .B(n644), .C(n195), .Y(n329) );
  NAND2X1 U265 ( .A(reg_array[38]), .B(n188), .Y(n195) );
  OAI21X1 U266 ( .A(n658), .B(n644), .C(n196), .Y(n330) );
  NAND2X1 U267 ( .A(reg_array[39]), .B(n188), .Y(n196) );
  OAI21X1 U268 ( .A(n657), .B(n644), .C(n197), .Y(n331) );
  NAND2X1 U269 ( .A(reg_array[40]), .B(n188), .Y(n197) );
  OAI21X1 U270 ( .A(n656), .B(n644), .C(n198), .Y(n332) );
  NAND2X1 U271 ( .A(reg_array[41]), .B(n188), .Y(n198) );
  OAI21X1 U272 ( .A(n655), .B(n644), .C(n199), .Y(n333) );
  NAND2X1 U273 ( .A(reg_array[42]), .B(n188), .Y(n199) );
  OAI21X1 U274 ( .A(n654), .B(n644), .C(n200), .Y(n334) );
  NAND2X1 U275 ( .A(reg_array[43]), .B(n188), .Y(n200) );
  OAI21X1 U276 ( .A(n653), .B(n188), .C(n201), .Y(n335) );
  NAND2X1 U277 ( .A(reg_array[44]), .B(n188), .Y(n201) );
  OAI21X1 U278 ( .A(n652), .B(n188), .C(n202), .Y(n336) );
  NAND2X1 U279 ( .A(reg_array[45]), .B(n188), .Y(n202) );
  OAI21X1 U280 ( .A(n651), .B(n188), .C(n203), .Y(n337) );
  NAND2X1 U281 ( .A(reg_array[46]), .B(n644), .Y(n203) );
  OAI21X1 U282 ( .A(n650), .B(n188), .C(n204), .Y(n338) );
  NAND2X1 U283 ( .A(reg_array[47]), .B(n644), .Y(n204) );
  NAND3X1 U284 ( .A(n170), .B(n668), .C(reg_write_dest[1]), .Y(n188) );
  OAI21X1 U285 ( .A(n665), .B(n642), .C(n206), .Y(n339) );
  NAND2X1 U286 ( .A(reg_array[48]), .B(n642), .Y(n206) );
  OAI21X1 U287 ( .A(n664), .B(n642), .C(n207), .Y(n340) );
  NAND2X1 U288 ( .A(reg_array[49]), .B(n642), .Y(n207) );
  OAI21X1 U289 ( .A(n663), .B(n642), .C(n208), .Y(n341) );
  NAND2X1 U290 ( .A(reg_array[50]), .B(n205), .Y(n208) );
  OAI21X1 U291 ( .A(n662), .B(n642), .C(n209), .Y(n342) );
  NAND2X1 U292 ( .A(reg_array[51]), .B(n205), .Y(n209) );
  OAI21X1 U293 ( .A(n661), .B(n642), .C(n210), .Y(n343) );
  NAND2X1 U294 ( .A(reg_array[52]), .B(n205), .Y(n210) );
  OAI21X1 U295 ( .A(n660), .B(n642), .C(n211), .Y(n344) );
  NAND2X1 U296 ( .A(reg_array[53]), .B(n205), .Y(n211) );
  OAI21X1 U297 ( .A(n659), .B(n642), .C(n212), .Y(n345) );
  NAND2X1 U298 ( .A(reg_array[54]), .B(n205), .Y(n212) );
  OAI21X1 U299 ( .A(n658), .B(n642), .C(n213), .Y(n346) );
  NAND2X1 U300 ( .A(reg_array[55]), .B(n205), .Y(n213) );
  OAI21X1 U301 ( .A(n657), .B(n642), .C(n214), .Y(n347) );
  NAND2X1 U302 ( .A(reg_array[56]), .B(n205), .Y(n214) );
  OAI21X1 U303 ( .A(n656), .B(n642), .C(n215), .Y(n348) );
  NAND2X1 U304 ( .A(reg_array[57]), .B(n205), .Y(n215) );
  OAI21X1 U305 ( .A(n655), .B(n642), .C(n216), .Y(n349) );
  NAND2X1 U306 ( .A(reg_array[58]), .B(n205), .Y(n216) );
  OAI21X1 U307 ( .A(n654), .B(n642), .C(n217), .Y(n350) );
  NAND2X1 U308 ( .A(reg_array[59]), .B(n205), .Y(n217) );
  OAI21X1 U309 ( .A(n653), .B(n205), .C(n218), .Y(n351) );
  NAND2X1 U310 ( .A(reg_array[60]), .B(n205), .Y(n218) );
  OAI21X1 U311 ( .A(n652), .B(n205), .C(n219), .Y(n352) );
  NAND2X1 U312 ( .A(reg_array[61]), .B(n205), .Y(n219) );
  OAI21X1 U313 ( .A(n651), .B(n205), .C(n220), .Y(n353) );
  NAND2X1 U314 ( .A(reg_array[62]), .B(n642), .Y(n220) );
  OAI21X1 U315 ( .A(n650), .B(n205), .C(n221), .Y(n354) );
  NAND2X1 U316 ( .A(reg_array[63]), .B(n642), .Y(n221) );
  NAND3X1 U317 ( .A(reg_write_dest[0]), .B(n170), .C(reg_write_dest[1]), .Y(
        n205) );
  NOR2X1 U318 ( .A(n666), .B(reg_write_dest[2]), .Y(n170) );
  OAI21X1 U319 ( .A(n665), .B(n640), .C(n223), .Y(n355) );
  NAND2X1 U320 ( .A(reg_array[64]), .B(n640), .Y(n223) );
  OAI21X1 U321 ( .A(n664), .B(n640), .C(n224), .Y(n356) );
  NAND2X1 U322 ( .A(reg_array[65]), .B(n640), .Y(n224) );
  OAI21X1 U323 ( .A(n663), .B(n640), .C(n225), .Y(n357) );
  NAND2X1 U324 ( .A(reg_array[66]), .B(n222), .Y(n225) );
  OAI21X1 U325 ( .A(n662), .B(n640), .C(n226), .Y(n358) );
  NAND2X1 U326 ( .A(reg_array[67]), .B(n222), .Y(n226) );
  OAI21X1 U327 ( .A(n661), .B(n640), .C(n227), .Y(n359) );
  NAND2X1 U328 ( .A(reg_array[68]), .B(n222), .Y(n227) );
  OAI21X1 U329 ( .A(n660), .B(n640), .C(n228), .Y(n360) );
  NAND2X1 U330 ( .A(reg_array[69]), .B(n222), .Y(n228) );
  OAI21X1 U331 ( .A(n659), .B(n640), .C(n229), .Y(n361) );
  NAND2X1 U332 ( .A(reg_array[70]), .B(n222), .Y(n229) );
  OAI21X1 U333 ( .A(n658), .B(n640), .C(n230), .Y(n362) );
  NAND2X1 U334 ( .A(reg_array[71]), .B(n222), .Y(n230) );
  OAI21X1 U335 ( .A(n657), .B(n640), .C(n231), .Y(n363) );
  NAND2X1 U336 ( .A(reg_array[72]), .B(n222), .Y(n231) );
  OAI21X1 U337 ( .A(n656), .B(n640), .C(n232), .Y(n364) );
  NAND2X1 U338 ( .A(reg_array[73]), .B(n222), .Y(n232) );
  OAI21X1 U339 ( .A(n655), .B(n640), .C(n233), .Y(n365) );
  NAND2X1 U340 ( .A(reg_array[74]), .B(n222), .Y(n233) );
  OAI21X1 U341 ( .A(n654), .B(n640), .C(n234), .Y(n366) );
  NAND2X1 U342 ( .A(reg_array[75]), .B(n222), .Y(n234) );
  OAI21X1 U343 ( .A(n653), .B(n222), .C(n235), .Y(n367) );
  NAND2X1 U344 ( .A(reg_array[76]), .B(n222), .Y(n235) );
  OAI21X1 U345 ( .A(n652), .B(n222), .C(n236), .Y(n368) );
  NAND2X1 U346 ( .A(reg_array[77]), .B(n222), .Y(n236) );
  OAI21X1 U347 ( .A(n651), .B(n222), .C(n237), .Y(n369) );
  NAND2X1 U348 ( .A(reg_array[78]), .B(n640), .Y(n237) );
  OAI21X1 U349 ( .A(n650), .B(n222), .C(n238), .Y(n370) );
  NAND2X1 U350 ( .A(reg_array[79]), .B(n640), .Y(n238) );
  NAND3X1 U351 ( .A(n668), .B(n667), .C(n239), .Y(n222) );
  OAI21X1 U352 ( .A(n665), .B(n638), .C(n241), .Y(n371) );
  NAND2X1 U353 ( .A(reg_array[80]), .B(n638), .Y(n241) );
  OAI21X1 U354 ( .A(n664), .B(n638), .C(n242), .Y(n372) );
  NAND2X1 U355 ( .A(reg_array[81]), .B(n638), .Y(n242) );
  OAI21X1 U356 ( .A(n663), .B(n638), .C(n243), .Y(n373) );
  NAND2X1 U357 ( .A(reg_array[82]), .B(n240), .Y(n243) );
  OAI21X1 U358 ( .A(n662), .B(n638), .C(n244), .Y(n374) );
  NAND2X1 U359 ( .A(reg_array[83]), .B(n240), .Y(n244) );
  OAI21X1 U360 ( .A(n661), .B(n638), .C(n245), .Y(n375) );
  NAND2X1 U361 ( .A(reg_array[84]), .B(n240), .Y(n245) );
  OAI21X1 U362 ( .A(n660), .B(n638), .C(n246), .Y(n376) );
  NAND2X1 U363 ( .A(reg_array[85]), .B(n240), .Y(n246) );
  OAI21X1 U364 ( .A(n659), .B(n638), .C(n247), .Y(n377) );
  NAND2X1 U365 ( .A(reg_array[86]), .B(n240), .Y(n247) );
  OAI21X1 U366 ( .A(n658), .B(n638), .C(n248), .Y(n378) );
  NAND2X1 U367 ( .A(reg_array[87]), .B(n240), .Y(n248) );
  OAI21X1 U368 ( .A(n657), .B(n638), .C(n249), .Y(n379) );
  NAND2X1 U369 ( .A(reg_array[88]), .B(n240), .Y(n249) );
  OAI21X1 U370 ( .A(n656), .B(n638), .C(n250), .Y(n380) );
  NAND2X1 U371 ( .A(reg_array[89]), .B(n240), .Y(n250) );
  OAI21X1 U372 ( .A(n655), .B(n638), .C(n251), .Y(n381) );
  NAND2X1 U373 ( .A(reg_array[90]), .B(n240), .Y(n251) );
  OAI21X1 U374 ( .A(n654), .B(n638), .C(n252), .Y(n382) );
  NAND2X1 U375 ( .A(reg_array[91]), .B(n240), .Y(n252) );
  OAI21X1 U376 ( .A(n653), .B(n240), .C(n253), .Y(n383) );
  NAND2X1 U377 ( .A(reg_array[92]), .B(n240), .Y(n253) );
  OAI21X1 U378 ( .A(n652), .B(n240), .C(n254), .Y(n384) );
  NAND2X1 U379 ( .A(reg_array[93]), .B(n240), .Y(n254) );
  OAI21X1 U380 ( .A(n651), .B(n240), .C(n255), .Y(n385) );
  NAND2X1 U381 ( .A(reg_array[94]), .B(n638), .Y(n255) );
  OAI21X1 U382 ( .A(n650), .B(n240), .C(n256), .Y(n386) );
  NAND2X1 U383 ( .A(reg_array[95]), .B(n638), .Y(n256) );
  NAND3X1 U384 ( .A(reg_write_dest[0]), .B(n667), .C(n239), .Y(n240) );
  OAI21X1 U385 ( .A(n665), .B(n636), .C(n258), .Y(n387) );
  NAND2X1 U386 ( .A(reg_array[96]), .B(n636), .Y(n258) );
  OAI21X1 U387 ( .A(n664), .B(n636), .C(n259), .Y(n388) );
  NAND2X1 U388 ( .A(reg_array[97]), .B(n636), .Y(n259) );
  OAI21X1 U389 ( .A(n663), .B(n636), .C(n260), .Y(n389) );
  NAND2X1 U390 ( .A(reg_array[98]), .B(n257), .Y(n260) );
  OAI21X1 U391 ( .A(n662), .B(n636), .C(n261), .Y(n390) );
  NAND2X1 U392 ( .A(reg_array[99]), .B(n257), .Y(n261) );
  OAI21X1 U393 ( .A(n661), .B(n636), .C(n262), .Y(n391) );
  NAND2X1 U394 ( .A(reg_array[100]), .B(n257), .Y(n262) );
  OAI21X1 U395 ( .A(n660), .B(n636), .C(n263), .Y(n392) );
  NAND2X1 U396 ( .A(reg_array[101]), .B(n257), .Y(n263) );
  OAI21X1 U397 ( .A(n659), .B(n636), .C(n264), .Y(n393) );
  NAND2X1 U398 ( .A(reg_array[102]), .B(n257), .Y(n264) );
  OAI21X1 U399 ( .A(n658), .B(n636), .C(n265), .Y(n394) );
  NAND2X1 U400 ( .A(reg_array[103]), .B(n257), .Y(n265) );
  OAI21X1 U401 ( .A(n657), .B(n636), .C(n266), .Y(n395) );
  NAND2X1 U402 ( .A(reg_array[104]), .B(n257), .Y(n266) );
  OAI21X1 U403 ( .A(n656), .B(n636), .C(n267), .Y(n396) );
  NAND2X1 U404 ( .A(reg_array[105]), .B(n257), .Y(n267) );
  OAI21X1 U405 ( .A(n655), .B(n636), .C(n268), .Y(n397) );
  NAND2X1 U406 ( .A(reg_array[106]), .B(n257), .Y(n268) );
  OAI21X1 U407 ( .A(n654), .B(n636), .C(n269), .Y(n398) );
  NAND2X1 U408 ( .A(reg_array[107]), .B(n257), .Y(n269) );
  OAI21X1 U409 ( .A(n653), .B(n257), .C(n270), .Y(n399) );
  NAND2X1 U410 ( .A(reg_array[108]), .B(n257), .Y(n270) );
  OAI21X1 U411 ( .A(n652), .B(n257), .C(n271), .Y(n400) );
  NAND2X1 U412 ( .A(reg_array[109]), .B(n257), .Y(n271) );
  OAI21X1 U413 ( .A(n651), .B(n257), .C(n272), .Y(n401) );
  NAND2X1 U414 ( .A(reg_array[110]), .B(n636), .Y(n272) );
  OAI21X1 U415 ( .A(n650), .B(n257), .C(n273), .Y(n402) );
  NAND2X1 U416 ( .A(reg_array[111]), .B(n636), .Y(n273) );
  NAND3X1 U417 ( .A(reg_write_dest[1]), .B(n668), .C(n239), .Y(n257) );
  OAI21X1 U418 ( .A(n665), .B(n634), .C(n275), .Y(n403) );
  NAND2X1 U419 ( .A(reg_array[112]), .B(n634), .Y(n275) );
  OAI21X1 U420 ( .A(n664), .B(n634), .C(n276), .Y(n404) );
  NAND2X1 U421 ( .A(reg_array[113]), .B(n634), .Y(n276) );
  OAI21X1 U422 ( .A(n663), .B(n634), .C(n277), .Y(n405) );
  NAND2X1 U423 ( .A(reg_array[114]), .B(n274), .Y(n277) );
  OAI21X1 U424 ( .A(n662), .B(n634), .C(n278), .Y(n406) );
  NAND2X1 U425 ( .A(reg_array[115]), .B(n274), .Y(n278) );
  OAI21X1 U426 ( .A(n661), .B(n634), .C(n279), .Y(n407) );
  NAND2X1 U427 ( .A(reg_array[116]), .B(n274), .Y(n279) );
  OAI21X1 U428 ( .A(n660), .B(n634), .C(n280), .Y(n408) );
  NAND2X1 U429 ( .A(reg_array[117]), .B(n274), .Y(n280) );
  OAI21X1 U430 ( .A(n659), .B(n634), .C(n281), .Y(n409) );
  NAND2X1 U431 ( .A(reg_array[118]), .B(n274), .Y(n281) );
  OAI21X1 U432 ( .A(n658), .B(n634), .C(n282), .Y(n410) );
  NAND2X1 U433 ( .A(reg_array[119]), .B(n274), .Y(n282) );
  OAI21X1 U434 ( .A(n657), .B(n634), .C(n283), .Y(n411) );
  NAND2X1 U435 ( .A(reg_array[120]), .B(n274), .Y(n283) );
  OAI21X1 U436 ( .A(n656), .B(n634), .C(n284), .Y(n412) );
  NAND2X1 U437 ( .A(reg_array[121]), .B(n274), .Y(n284) );
  OAI21X1 U438 ( .A(n655), .B(n634), .C(n285), .Y(n413) );
  NAND2X1 U439 ( .A(reg_array[122]), .B(n274), .Y(n285) );
  OAI21X1 U440 ( .A(n654), .B(n634), .C(n286), .Y(n414) );
  NAND2X1 U441 ( .A(reg_array[123]), .B(n274), .Y(n286) );
  OAI21X1 U442 ( .A(n653), .B(n274), .C(n287), .Y(n415) );
  NAND2X1 U443 ( .A(reg_array[124]), .B(n274), .Y(n287) );
  OAI21X1 U444 ( .A(n652), .B(n274), .C(n288), .Y(n416) );
  NAND2X1 U445 ( .A(reg_array[125]), .B(n274), .Y(n288) );
  OAI21X1 U446 ( .A(n651), .B(n274), .C(n289), .Y(n417) );
  NAND2X1 U447 ( .A(reg_array[126]), .B(n634), .Y(n289) );
  OAI21X1 U448 ( .A(n650), .B(n274), .C(n290), .Y(n418) );
  NAND2X1 U449 ( .A(reg_array[127]), .B(n634), .Y(n290) );
  NAND3X1 U450 ( .A(reg_write_dest[1]), .B(reg_write_dest[0]), .C(n239), .Y(
        n274) );
  AND2X1 U451 ( .A(reg_write_dest[2]), .B(reg_write_en), .Y(n239) );
  BUFX2 U129 ( .A(reg_read_addr_1[1]), .Y(n128) );
  INVX2 U131 ( .A(n624), .Y(n625) );
  INVX2 U132 ( .A(n641), .Y(n640) );
  INVX2 U133 ( .A(n649), .Y(n648) );
  BUFX2 U134 ( .A(n633), .Y(n632) );
  BUFX2 U135 ( .A(n630), .Y(n633) );
  BUFX2 U136 ( .A(reg_read_addr_2[0]), .Y(n627) );
  INVX2 U137 ( .A(reg_read_addr_2[1]), .Y(n624) );
  INVX2 U138 ( .A(n629), .Y(n628) );
  BUFX2 U139 ( .A(reg_read_addr_2[0]), .Y(n626) );
  INVX2 U140 ( .A(n153), .Y(n649) );
  INVX2 U141 ( .A(n222), .Y(n641) );
  INVX2 U142 ( .A(n647), .Y(n646) );
  INVX2 U143 ( .A(n645), .Y(n644) );
  INVX2 U144 ( .A(n643), .Y(n642) );
  INVX2 U145 ( .A(n639), .Y(n638) );
  INVX2 U146 ( .A(n637), .Y(n636) );
  INVX2 U147 ( .A(n635), .Y(n634) );
  BUFX2 U148 ( .A(n671), .Y(n630) );
  BUFX2 U149 ( .A(n671), .Y(n631) );
  BUFX2 U150 ( .A(reg_read_addr_1[0]), .Y(n511) );
  BUFX2 U151 ( .A(reg_read_addr_1[0]), .Y(n510) );
  INVX2 U452 ( .A(n151), .Y(n669) );
  INVX2 U453 ( .A(reg_read_addr_2[2]), .Y(n629) );
  INVX2 U454 ( .A(n171), .Y(n647) );
  INVX2 U455 ( .A(n188), .Y(n645) );
  INVX2 U456 ( .A(n205), .Y(n643) );
  INVX2 U457 ( .A(n240), .Y(n639) );
  INVX2 U458 ( .A(n257), .Y(n637) );
  INVX2 U459 ( .A(n274), .Y(n635) );
  INVX2 U460 ( .A(n152), .Y(n670) );
  MUX2X1 U461 ( .B(n131), .A(n132), .S(n128), .Y(n130) );
  MUX2X1 U462 ( .B(n134), .A(n135), .S(n128), .Y(n133) );
  MUX2X1 U463 ( .B(n137), .A(n138), .S(n128), .Y(n136) );
  MUX2X1 U464 ( .B(n140), .A(n141), .S(n128), .Y(n139) );
  MUX2X1 U465 ( .B(n143), .A(n144), .S(n128), .Y(n142) );
  MUX2X1 U466 ( .B(n146), .A(n147), .S(n128), .Y(n145) );
  MUX2X1 U467 ( .B(n149), .A(n150), .S(n128), .Y(n148) );
  MUX2X1 U468 ( .B(n420), .A(n421), .S(n128), .Y(n419) );
  MUX2X1 U469 ( .B(n423), .A(n424), .S(n128), .Y(n422) );
  MUX2X1 U470 ( .B(n426), .A(n427), .S(n128), .Y(n425) );
  MUX2X1 U471 ( .B(n429), .A(n430), .S(n128), .Y(n428) );
  MUX2X1 U472 ( .B(n432), .A(n433), .S(n128), .Y(n431) );
  MUX2X1 U473 ( .B(n435), .A(n436), .S(n128), .Y(n434) );
  MUX2X1 U474 ( .B(n438), .A(n439), .S(n128), .Y(n437) );
  MUX2X1 U475 ( .B(n441), .A(n442), .S(n128), .Y(n440) );
  MUX2X1 U476 ( .B(n444), .A(n445), .S(n128), .Y(n443) );
  MUX2X1 U477 ( .B(n447), .A(n448), .S(n128), .Y(n446) );
  MUX2X1 U478 ( .B(n450), .A(n451), .S(n128), .Y(n449) );
  MUX2X1 U479 ( .B(n453), .A(n454), .S(n128), .Y(n452) );
  MUX2X1 U480 ( .B(n456), .A(n457), .S(n128), .Y(n455) );
  MUX2X1 U481 ( .B(n459), .A(n460), .S(n128), .Y(n458) );
  MUX2X1 U482 ( .B(n462), .A(n463), .S(n128), .Y(n461) );
  MUX2X1 U483 ( .B(n465), .A(n466), .S(n128), .Y(n464) );
  MUX2X1 U484 ( .B(n468), .A(n469), .S(n128), .Y(n467) );
  MUX2X1 U485 ( .B(n471), .A(n472), .S(n128), .Y(n470) );
  MUX2X1 U486 ( .B(n474), .A(n475), .S(n128), .Y(n473) );
  MUX2X1 U487 ( .B(n477), .A(n478), .S(n128), .Y(n476) );
  MUX2X1 U488 ( .B(n480), .A(n481), .S(n128), .Y(n479) );
  MUX2X1 U489 ( .B(n483), .A(n484), .S(n128), .Y(n482) );
  MUX2X1 U490 ( .B(n486), .A(n487), .S(n128), .Y(n485) );
  MUX2X1 U491 ( .B(n489), .A(n490), .S(n128), .Y(n488) );
  MUX2X1 U492 ( .B(n492), .A(n493), .S(n128), .Y(n491) );
  MUX2X1 U493 ( .B(reg_array[96]), .A(reg_array[112]), .S(n510), .Y(n132) );
  MUX2X1 U494 ( .B(reg_array[64]), .A(reg_array[80]), .S(n510), .Y(n131) );
  MUX2X1 U495 ( .B(reg_array[32]), .A(reg_array[48]), .S(reg_read_addr_1[0]), 
        .Y(n135) );
  MUX2X1 U496 ( .B(reg_array[0]), .A(reg_array[16]), .S(reg_read_addr_1[0]), 
        .Y(n134) );
  MUX2X1 U497 ( .B(n133), .A(n130), .S(reg_read_addr_1[2]), .Y(n494) );
  INVX2 U498 ( .A(n494), .Y(N44) );
  MUX2X1 U499 ( .B(reg_array[97]), .A(reg_array[113]), .S(reg_read_addr_1[0]), 
        .Y(n138) );
  MUX2X1 U500 ( .B(reg_array[65]), .A(reg_array[81]), .S(reg_read_addr_1[0]), 
        .Y(n137) );
  MUX2X1 U501 ( .B(reg_array[33]), .A(reg_array[49]), .S(reg_read_addr_1[0]), 
        .Y(n141) );
  MUX2X1 U502 ( .B(reg_array[1]), .A(reg_array[17]), .S(reg_read_addr_1[0]), 
        .Y(n140) );
  MUX2X1 U503 ( .B(n139), .A(n136), .S(reg_read_addr_1[2]), .Y(n495) );
  INVX2 U504 ( .A(n495), .Y(N43) );
  MUX2X1 U505 ( .B(reg_array[98]), .A(reg_array[114]), .S(n511), .Y(n144) );
  MUX2X1 U506 ( .B(reg_array[66]), .A(reg_array[82]), .S(n510), .Y(n143) );
  MUX2X1 U507 ( .B(reg_array[34]), .A(reg_array[50]), .S(n511), .Y(n147) );
  MUX2X1 U508 ( .B(reg_array[2]), .A(reg_array[18]), .S(n510), .Y(n146) );
  MUX2X1 U509 ( .B(n145), .A(n142), .S(reg_read_addr_1[2]), .Y(n496) );
  INVX2 U510 ( .A(n496), .Y(N42) );
  MUX2X1 U511 ( .B(reg_array[99]), .A(reg_array[115]), .S(n511), .Y(n150) );
  MUX2X1 U512 ( .B(reg_array[67]), .A(reg_array[83]), .S(reg_read_addr_1[0]), 
        .Y(n149) );
  MUX2X1 U513 ( .B(reg_array[35]), .A(reg_array[51]), .S(reg_read_addr_1[0]), 
        .Y(n421) );
  MUX2X1 U514 ( .B(reg_array[3]), .A(reg_array[19]), .S(n511), .Y(n420) );
  MUX2X1 U515 ( .B(n419), .A(n148), .S(reg_read_addr_1[2]), .Y(n497) );
  INVX2 U516 ( .A(n497), .Y(N41) );
  MUX2X1 U517 ( .B(reg_array[100]), .A(reg_array[116]), .S(n510), .Y(n424) );
  MUX2X1 U518 ( .B(reg_array[68]), .A(reg_array[84]), .S(n510), .Y(n423) );
  MUX2X1 U519 ( .B(reg_array[36]), .A(reg_array[52]), .S(n510), .Y(n427) );
  MUX2X1 U520 ( .B(reg_array[4]), .A(reg_array[20]), .S(n510), .Y(n426) );
  MUX2X1 U521 ( .B(n425), .A(n422), .S(reg_read_addr_1[2]), .Y(n498) );
  INVX2 U522 ( .A(n498), .Y(N40) );
  MUX2X1 U523 ( .B(reg_array[101]), .A(reg_array[117]), .S(n510), .Y(n430) );
  MUX2X1 U524 ( .B(reg_array[69]), .A(reg_array[85]), .S(n510), .Y(n429) );
  MUX2X1 U525 ( .B(reg_array[37]), .A(reg_array[53]), .S(n510), .Y(n433) );
  MUX2X1 U526 ( .B(reg_array[5]), .A(reg_array[21]), .S(n510), .Y(n432) );
  MUX2X1 U527 ( .B(n431), .A(n428), .S(reg_read_addr_1[2]), .Y(n499) );
  INVX2 U528 ( .A(n499), .Y(N39) );
  MUX2X1 U529 ( .B(reg_array[102]), .A(reg_array[118]), .S(n510), .Y(n436) );
  MUX2X1 U530 ( .B(reg_array[70]), .A(reg_array[86]), .S(n510), .Y(n435) );
  MUX2X1 U531 ( .B(reg_array[38]), .A(reg_array[54]), .S(n510), .Y(n439) );
  MUX2X1 U532 ( .B(reg_array[6]), .A(reg_array[22]), .S(n510), .Y(n438) );
  MUX2X1 U533 ( .B(n437), .A(n434), .S(reg_read_addr_1[2]), .Y(n500) );
  INVX2 U534 ( .A(n500), .Y(N38) );
  MUX2X1 U535 ( .B(reg_array[103]), .A(reg_array[119]), .S(n511), .Y(n442) );
  MUX2X1 U536 ( .B(reg_array[71]), .A(reg_array[87]), .S(n511), .Y(n441) );
  MUX2X1 U537 ( .B(reg_array[39]), .A(reg_array[55]), .S(n511), .Y(n445) );
  MUX2X1 U538 ( .B(reg_array[7]), .A(reg_array[23]), .S(n511), .Y(n444) );
  MUX2X1 U539 ( .B(n443), .A(n440), .S(reg_read_addr_1[2]), .Y(n501) );
  INVX2 U540 ( .A(n501), .Y(N37) );
  MUX2X1 U541 ( .B(reg_array[104]), .A(reg_array[120]), .S(n511), .Y(n448) );
  MUX2X1 U542 ( .B(reg_array[72]), .A(reg_array[88]), .S(n511), .Y(n447) );
  MUX2X1 U543 ( .B(reg_array[40]), .A(reg_array[56]), .S(n511), .Y(n451) );
  MUX2X1 U544 ( .B(reg_array[8]), .A(reg_array[24]), .S(n511), .Y(n450) );
  MUX2X1 U545 ( .B(n449), .A(n446), .S(reg_read_addr_1[2]), .Y(n502) );
  INVX2 U546 ( .A(n502), .Y(N36) );
  MUX2X1 U547 ( .B(reg_array[105]), .A(reg_array[121]), .S(n511), .Y(n454) );
  MUX2X1 U548 ( .B(reg_array[73]), .A(reg_array[89]), .S(n511), .Y(n453) );
  MUX2X1 U549 ( .B(reg_array[41]), .A(reg_array[57]), .S(n511), .Y(n457) );
  MUX2X1 U550 ( .B(reg_array[9]), .A(reg_array[25]), .S(n511), .Y(n456) );
  MUX2X1 U551 ( .B(n455), .A(n452), .S(reg_read_addr_1[2]), .Y(n503) );
  INVX2 U552 ( .A(n503), .Y(N35) );
  MUX2X1 U553 ( .B(reg_array[106]), .A(reg_array[122]), .S(reg_read_addr_1[0]), 
        .Y(n460) );
  MUX2X1 U554 ( .B(reg_array[74]), .A(reg_array[90]), .S(n510), .Y(n459) );
  MUX2X1 U555 ( .B(reg_array[42]), .A(reg_array[58]), .S(reg_read_addr_1[0]), 
        .Y(n463) );
  MUX2X1 U556 ( .B(reg_array[10]), .A(reg_array[26]), .S(n511), .Y(n462) );
  MUX2X1 U557 ( .B(n461), .A(n458), .S(reg_read_addr_1[2]), .Y(n504) );
  INVX2 U558 ( .A(n504), .Y(N34) );
  MUX2X1 U559 ( .B(reg_array[107]), .A(reg_array[123]), .S(reg_read_addr_1[0]), 
        .Y(n466) );
  MUX2X1 U560 ( .B(reg_array[75]), .A(reg_array[91]), .S(reg_read_addr_1[0]), 
        .Y(n465) );
  MUX2X1 U561 ( .B(reg_array[43]), .A(reg_array[59]), .S(reg_read_addr_1[0]), 
        .Y(n469) );
  MUX2X1 U562 ( .B(reg_array[11]), .A(reg_array[27]), .S(reg_read_addr_1[0]), 
        .Y(n468) );
  MUX2X1 U563 ( .B(n467), .A(n464), .S(reg_read_addr_1[2]), .Y(n505) );
  INVX2 U564 ( .A(n505), .Y(N33) );
  MUX2X1 U565 ( .B(reg_array[108]), .A(reg_array[124]), .S(n511), .Y(n472) );
  MUX2X1 U566 ( .B(reg_array[76]), .A(reg_array[92]), .S(n510), .Y(n471) );
  MUX2X1 U567 ( .B(reg_array[44]), .A(reg_array[60]), .S(n510), .Y(n475) );
  MUX2X1 U568 ( .B(reg_array[12]), .A(reg_array[28]), .S(n511), .Y(n474) );
  MUX2X1 U569 ( .B(n473), .A(n470), .S(reg_read_addr_1[2]), .Y(n506) );
  INVX2 U570 ( .A(n506), .Y(N32) );
  MUX2X1 U571 ( .B(reg_array[109]), .A(reg_array[125]), .S(n511), .Y(n478) );
  MUX2X1 U572 ( .B(reg_array[77]), .A(reg_array[93]), .S(n511), .Y(n477) );
  MUX2X1 U573 ( .B(reg_array[45]), .A(reg_array[61]), .S(n510), .Y(n481) );
  MUX2X1 U574 ( .B(reg_array[13]), .A(reg_array[29]), .S(n510), .Y(n480) );
  MUX2X1 U575 ( .B(n479), .A(n476), .S(reg_read_addr_1[2]), .Y(n507) );
  INVX2 U576 ( .A(n507), .Y(N31) );
  MUX2X1 U577 ( .B(reg_array[110]), .A(reg_array[126]), .S(n511), .Y(n484) );
  MUX2X1 U578 ( .B(reg_array[78]), .A(reg_array[94]), .S(n511), .Y(n483) );
  MUX2X1 U579 ( .B(reg_array[46]), .A(reg_array[62]), .S(n510), .Y(n487) );
  MUX2X1 U580 ( .B(reg_array[14]), .A(reg_array[30]), .S(n510), .Y(n486) );
  MUX2X1 U581 ( .B(n485), .A(n482), .S(reg_read_addr_1[2]), .Y(n508) );
  INVX2 U582 ( .A(n508), .Y(N30) );
  MUX2X1 U583 ( .B(reg_array[111]), .A(reg_array[127]), .S(n511), .Y(n490) );
  MUX2X1 U584 ( .B(reg_array[79]), .A(reg_array[95]), .S(n511), .Y(n489) );
  MUX2X1 U585 ( .B(reg_array[47]), .A(reg_array[63]), .S(n510), .Y(n493) );
  MUX2X1 U586 ( .B(reg_array[15]), .A(reg_array[31]), .S(n510), .Y(n492) );
  MUX2X1 U587 ( .B(n491), .A(n488), .S(reg_read_addr_1[2]), .Y(n509) );
  INVX2 U588 ( .A(n509), .Y(N29) );
  MUX2X1 U589 ( .B(n513), .A(n514), .S(reg_read_addr_2[1]), .Y(n512) );
  MUX2X1 U590 ( .B(n516), .A(n517), .S(n625), .Y(n515) );
  MUX2X1 U591 ( .B(n519), .A(n520), .S(reg_read_addr_2[1]), .Y(n518) );
  MUX2X1 U592 ( .B(n522), .A(n523), .S(n625), .Y(n521) );
  MUX2X1 U593 ( .B(n525), .A(n526), .S(reg_read_addr_2[1]), .Y(n524) );
  MUX2X1 U594 ( .B(n528), .A(n529), .S(n625), .Y(n527) );
  MUX2X1 U595 ( .B(n531), .A(n532), .S(reg_read_addr_2[1]), .Y(n530) );
  MUX2X1 U596 ( .B(n534), .A(n535), .S(reg_read_addr_2[1]), .Y(n533) );
  MUX2X1 U597 ( .B(n537), .A(n538), .S(n625), .Y(n536) );
  MUX2X1 U598 ( .B(n540), .A(n541), .S(reg_read_addr_2[1]), .Y(n539) );
  MUX2X1 U599 ( .B(n543), .A(n544), .S(reg_read_addr_2[1]), .Y(n542) );
  MUX2X1 U600 ( .B(n546), .A(n547), .S(reg_read_addr_2[1]), .Y(n545) );
  MUX2X1 U601 ( .B(n549), .A(n550), .S(n625), .Y(n548) );
  MUX2X1 U602 ( .B(n552), .A(n553), .S(n625), .Y(n551) );
  MUX2X1 U603 ( .B(n555), .A(n556), .S(n625), .Y(n554) );
  MUX2X1 U604 ( .B(n558), .A(n559), .S(n625), .Y(n557) );
  MUX2X1 U605 ( .B(n561), .A(n562), .S(n625), .Y(n560) );
  MUX2X1 U606 ( .B(n564), .A(n565), .S(n625), .Y(n563) );
  MUX2X1 U607 ( .B(n567), .A(n568), .S(n625), .Y(n566) );
  MUX2X1 U608 ( .B(n570), .A(n571), .S(n625), .Y(n569) );
  MUX2X1 U609 ( .B(n573), .A(n574), .S(n625), .Y(n572) );
  MUX2X1 U610 ( .B(n576), .A(n577), .S(n625), .Y(n575) );
  MUX2X1 U611 ( .B(n579), .A(n580), .S(n625), .Y(n578) );
  MUX2X1 U612 ( .B(n582), .A(n583), .S(n625), .Y(n581) );
  MUX2X1 U613 ( .B(n585), .A(n586), .S(reg_read_addr_2[1]), .Y(n584) );
  MUX2X1 U614 ( .B(n588), .A(n589), .S(reg_read_addr_2[1]), .Y(n587) );
  MUX2X1 U615 ( .B(n591), .A(n592), .S(n625), .Y(n590) );
  MUX2X1 U616 ( .B(n594), .A(n595), .S(reg_read_addr_2[1]), .Y(n593) );
  MUX2X1 U617 ( .B(n597), .A(n598), .S(reg_read_addr_2[1]), .Y(n596) );
  MUX2X1 U618 ( .B(n600), .A(n601), .S(reg_read_addr_2[1]), .Y(n599) );
  MUX2X1 U619 ( .B(n603), .A(n604), .S(n625), .Y(n602) );
  MUX2X1 U620 ( .B(n606), .A(n607), .S(reg_read_addr_2[1]), .Y(n605) );
  MUX2X1 U621 ( .B(reg_array[96]), .A(reg_array[112]), .S(n626), .Y(n514) );
  MUX2X1 U622 ( .B(reg_array[64]), .A(reg_array[80]), .S(n626), .Y(n513) );
  MUX2X1 U623 ( .B(reg_array[32]), .A(reg_array[48]), .S(n626), .Y(n517) );
  MUX2X1 U624 ( .B(reg_array[0]), .A(reg_array[16]), .S(n626), .Y(n516) );
  MUX2X1 U625 ( .B(n515), .A(n512), .S(n628), .Y(n608) );
  INVX2 U626 ( .A(n608), .Y(N60) );
  MUX2X1 U627 ( .B(reg_array[97]), .A(reg_array[113]), .S(n626), .Y(n520) );
  MUX2X1 U628 ( .B(reg_array[65]), .A(reg_array[81]), .S(n627), .Y(n519) );
  MUX2X1 U629 ( .B(reg_array[33]), .A(reg_array[49]), .S(n626), .Y(n523) );
  MUX2X1 U630 ( .B(reg_array[1]), .A(reg_array[17]), .S(n627), .Y(n522) );
  MUX2X1 U631 ( .B(n521), .A(n518), .S(reg_read_addr_2[2]), .Y(n609) );
  INVX2 U632 ( .A(n609), .Y(N59) );
  MUX2X1 U633 ( .B(reg_array[98]), .A(reg_array[114]), .S(n627), .Y(n526) );
  MUX2X1 U634 ( .B(reg_array[66]), .A(reg_array[82]), .S(n626), .Y(n525) );
  MUX2X1 U635 ( .B(reg_array[34]), .A(reg_array[50]), .S(n627), .Y(n529) );
  MUX2X1 U636 ( .B(reg_array[2]), .A(reg_array[18]), .S(n626), .Y(n528) );
  MUX2X1 U637 ( .B(n527), .A(n524), .S(n628), .Y(n610) );
  INVX2 U638 ( .A(n610), .Y(N58) );
  MUX2X1 U639 ( .B(reg_array[99]), .A(reg_array[115]), .S(n626), .Y(n532) );
  MUX2X1 U640 ( .B(reg_array[67]), .A(reg_array[83]), .S(n626), .Y(n531) );
  MUX2X1 U641 ( .B(reg_array[35]), .A(reg_array[51]), .S(n626), .Y(n535) );
  MUX2X1 U642 ( .B(reg_array[3]), .A(reg_array[19]), .S(n627), .Y(n534) );
  MUX2X1 U643 ( .B(n533), .A(n530), .S(n628), .Y(n611) );
  INVX2 U644 ( .A(n611), .Y(N57) );
  MUX2X1 U645 ( .B(reg_array[100]), .A(reg_array[116]), .S(n626), .Y(n538) );
  MUX2X1 U646 ( .B(reg_array[68]), .A(reg_array[84]), .S(n627), .Y(n537) );
  MUX2X1 U647 ( .B(reg_array[36]), .A(reg_array[52]), .S(n627), .Y(n541) );
  MUX2X1 U648 ( .B(reg_array[4]), .A(reg_array[20]), .S(n627), .Y(n540) );
  MUX2X1 U649 ( .B(n539), .A(n536), .S(n628), .Y(n612) );
  INVX2 U650 ( .A(n612), .Y(N56) );
  MUX2X1 U651 ( .B(reg_array[101]), .A(reg_array[117]), .S(reg_read_addr_2[0]), 
        .Y(n544) );
  MUX2X1 U652 ( .B(reg_array[69]), .A(reg_array[85]), .S(n627), .Y(n543) );
  MUX2X1 U653 ( .B(reg_array[37]), .A(reg_array[53]), .S(reg_read_addr_2[0]), 
        .Y(n547) );
  MUX2X1 U654 ( .B(reg_array[5]), .A(reg_array[21]), .S(reg_read_addr_2[0]), 
        .Y(n546) );
  MUX2X1 U655 ( .B(n545), .A(n542), .S(reg_read_addr_2[2]), .Y(n613) );
  INVX2 U656 ( .A(n613), .Y(N55) );
  MUX2X1 U657 ( .B(reg_array[102]), .A(reg_array[118]), .S(reg_read_addr_2[0]), 
        .Y(n550) );
  MUX2X1 U658 ( .B(reg_array[70]), .A(reg_array[86]), .S(n626), .Y(n549) );
  MUX2X1 U659 ( .B(reg_array[38]), .A(reg_array[54]), .S(reg_read_addr_2[0]), 
        .Y(n553) );
  MUX2X1 U660 ( .B(reg_array[6]), .A(reg_array[22]), .S(reg_read_addr_2[0]), 
        .Y(n552) );
  MUX2X1 U661 ( .B(n551), .A(n548), .S(n628), .Y(n614) );
  INVX2 U662 ( .A(n614), .Y(N54) );
  MUX2X1 U663 ( .B(reg_array[103]), .A(reg_array[119]), .S(reg_read_addr_2[0]), 
        .Y(n556) );
  MUX2X1 U664 ( .B(reg_array[71]), .A(reg_array[87]), .S(reg_read_addr_2[0]), 
        .Y(n555) );
  MUX2X1 U665 ( .B(reg_array[39]), .A(reg_array[55]), .S(reg_read_addr_2[0]), 
        .Y(n559) );
  MUX2X1 U666 ( .B(reg_array[7]), .A(reg_array[23]), .S(n627), .Y(n558) );
  MUX2X1 U667 ( .B(n557), .A(n554), .S(reg_read_addr_2[2]), .Y(n615) );
  INVX2 U668 ( .A(n615), .Y(N53) );
  MUX2X1 U669 ( .B(reg_array[104]), .A(reg_array[120]), .S(n626), .Y(n562) );
  MUX2X1 U670 ( .B(reg_array[72]), .A(reg_array[88]), .S(reg_read_addr_2[0]), 
        .Y(n561) );
  MUX2X1 U671 ( .B(reg_array[40]), .A(reg_array[56]), .S(n627), .Y(n565) );
  MUX2X1 U672 ( .B(reg_array[8]), .A(reg_array[24]), .S(reg_read_addr_2[0]), 
        .Y(n564) );
  MUX2X1 U673 ( .B(n563), .A(n560), .S(n628), .Y(n616) );
  INVX2 U674 ( .A(n616), .Y(N52) );
  MUX2X1 U675 ( .B(reg_array[105]), .A(reg_array[121]), .S(n626), .Y(n568) );
  MUX2X1 U676 ( .B(reg_array[73]), .A(reg_array[89]), .S(reg_read_addr_2[0]), 
        .Y(n567) );
  MUX2X1 U677 ( .B(reg_array[41]), .A(reg_array[57]), .S(n626), .Y(n571) );
  MUX2X1 U678 ( .B(reg_array[9]), .A(reg_array[25]), .S(reg_read_addr_2[0]), 
        .Y(n570) );
  MUX2X1 U679 ( .B(n569), .A(n566), .S(reg_read_addr_2[2]), .Y(n617) );
  INVX2 U680 ( .A(n617), .Y(N51) );
  MUX2X1 U681 ( .B(reg_array[106]), .A(reg_array[122]), .S(n626), .Y(n574) );
  MUX2X1 U682 ( .B(reg_array[74]), .A(reg_array[90]), .S(n627), .Y(n573) );
  MUX2X1 U683 ( .B(reg_array[42]), .A(reg_array[58]), .S(n626), .Y(n577) );
  MUX2X1 U684 ( .B(reg_array[10]), .A(reg_array[26]), .S(n627), .Y(n576) );
  MUX2X1 U685 ( .B(n575), .A(n572), .S(n628), .Y(n618) );
  INVX2 U686 ( .A(n618), .Y(N50) );
  MUX2X1 U687 ( .B(reg_array[107]), .A(reg_array[123]), .S(n626), .Y(n580) );
  MUX2X1 U688 ( .B(reg_array[75]), .A(reg_array[91]), .S(n626), .Y(n579) );
  MUX2X1 U689 ( .B(reg_array[43]), .A(reg_array[59]), .S(n626), .Y(n583) );
  MUX2X1 U690 ( .B(reg_array[11]), .A(reg_array[27]), .S(n626), .Y(n582) );
  MUX2X1 U691 ( .B(n581), .A(n578), .S(reg_read_addr_2[2]), .Y(n619) );
  INVX2 U692 ( .A(n619), .Y(N49) );
  MUX2X1 U693 ( .B(reg_array[108]), .A(reg_array[124]), .S(n626), .Y(n586) );
  MUX2X1 U694 ( .B(reg_array[76]), .A(reg_array[92]), .S(reg_read_addr_2[0]), 
        .Y(n585) );
  MUX2X1 U695 ( .B(reg_array[44]), .A(reg_array[60]), .S(n626), .Y(n589) );
  MUX2X1 U696 ( .B(reg_array[12]), .A(reg_array[28]), .S(n626), .Y(n588) );
  MUX2X1 U697 ( .B(n587), .A(n584), .S(n628), .Y(n620) );
  INVX2 U698 ( .A(n620), .Y(N48) );
  MUX2X1 U699 ( .B(reg_array[109]), .A(reg_array[125]), .S(n627), .Y(n592) );
  MUX2X1 U700 ( .B(reg_array[77]), .A(reg_array[93]), .S(n627), .Y(n591) );
  MUX2X1 U701 ( .B(reg_array[45]), .A(reg_array[61]), .S(n627), .Y(n595) );
  MUX2X1 U702 ( .B(reg_array[13]), .A(reg_array[29]), .S(n627), .Y(n594) );
  MUX2X1 U703 ( .B(n593), .A(n590), .S(reg_read_addr_2[2]), .Y(n621) );
  INVX2 U704 ( .A(n621), .Y(N47) );
  MUX2X1 U705 ( .B(reg_array[110]), .A(reg_array[126]), .S(n627), .Y(n598) );
  MUX2X1 U706 ( .B(reg_array[78]), .A(reg_array[94]), .S(n627), .Y(n597) );
  MUX2X1 U707 ( .B(reg_array[46]), .A(reg_array[62]), .S(n627), .Y(n601) );
  MUX2X1 U708 ( .B(reg_array[14]), .A(reg_array[30]), .S(n627), .Y(n600) );
  MUX2X1 U709 ( .B(n599), .A(n596), .S(n628), .Y(n622) );
  INVX2 U710 ( .A(n622), .Y(N46) );
  MUX2X1 U711 ( .B(reg_array[111]), .A(reg_array[127]), .S(n627), .Y(n604) );
  MUX2X1 U712 ( .B(reg_array[79]), .A(reg_array[95]), .S(n627), .Y(n603) );
  MUX2X1 U713 ( .B(reg_array[47]), .A(reg_array[63]), .S(n627), .Y(n607) );
  MUX2X1 U714 ( .B(reg_array[15]), .A(reg_array[31]), .S(n627), .Y(n606) );
  MUX2X1 U715 ( .B(n605), .A(n602), .S(reg_read_addr_2[2]), .Y(n623) );
  INVX2 U716 ( .A(n623), .Y(N45) );
  INVX2 U717 ( .A(reg_write_data[15]), .Y(n650) );
  INVX2 U718 ( .A(reg_write_data[14]), .Y(n651) );
  INVX2 U719 ( .A(reg_write_data[13]), .Y(n652) );
  INVX2 U720 ( .A(reg_write_data[12]), .Y(n653) );
  INVX2 U721 ( .A(reg_write_data[11]), .Y(n654) );
  INVX2 U722 ( .A(reg_write_data[10]), .Y(n655) );
  INVX2 U723 ( .A(reg_write_data[9]), .Y(n656) );
  INVX2 U724 ( .A(reg_write_data[8]), .Y(n657) );
  INVX2 U725 ( .A(reg_write_data[7]), .Y(n658) );
  INVX2 U726 ( .A(reg_write_data[6]), .Y(n659) );
  INVX2 U727 ( .A(reg_write_data[5]), .Y(n660) );
  INVX2 U728 ( .A(reg_write_data[4]), .Y(n661) );
  INVX2 U729 ( .A(reg_write_data[3]), .Y(n662) );
  INVX2 U730 ( .A(reg_write_data[2]), .Y(n663) );
  INVX2 U731 ( .A(reg_write_data[1]), .Y(n664) );
  INVX2 U732 ( .A(reg_write_data[0]), .Y(n665) );
  INVX2 U733 ( .A(reg_write_en), .Y(n666) );
  INVX2 U734 ( .A(reg_write_dest[1]), .Y(n667) );
  INVX2 U735 ( .A(reg_write_dest[0]), .Y(n668) );
  INVX2 U736 ( .A(rst), .Y(n671) );
endmodule


module FSM ( clk, rst, pc );
  output [7:0] pc;
  input clk, rst;
  wire   instruction_fetch_en, branch_taken, baseline_en, reg_write_en, n1, n3,
         n4, SYNOPSYS_UNCONNECTED_1;
  wire   [5:0] branch_offset_imm;
  wire   [15:0] instruction;
  wire   [57:0] ID_pipeline_reg_out;
  wire   [2:0] reg_read_addr_1;
  wire   [2:0] reg_read_addr_2;
  wire   [15:0] reg_read_data_1;
  wire   [15:0] reg_read_data_2;
  wire   [38:0] EX_pipeline_reg_out;
  wire   [37:0] MEM_pipeline_reg_out;
  wire   [2:0] reg_write_dest;
  wire   [15:0] reg_write_data;

  IF_stage IF_stage_inst ( .clk(clk), .rst(n4), .instruction_fetch_en(
        instruction_fetch_en), .branch_offset_imm(branch_offset_imm), 
        .branch_taken(branch_taken), .pc(pc), .instruction({instruction[15:3], 
        SYNOPSYS_UNCONNECTED_1, instruction[1:0]}), .baseline_en(baseline_en)
         );
  ID_stage ID_stage_inst ( .clk(clk), .rst(n4), .baseline_en(baseline_en), 
        .pipeline_reg_out(ID_pipeline_reg_out), .instruction({
        instruction[15:3], 1'b0, instruction[1:0]}), .branch_offset_imm(
        branch_offset_imm), .branch_taken(branch_taken), .reg_read_addr_1(
        reg_read_addr_1), .reg_read_addr_2(reg_read_addr_2), .reg_read_data_1(
        reg_read_data_1), .reg_read_data_2(reg_read_data_2) );
  EX_stage EX_stage_inst ( .clk(clk), .rst(n4), .pipeline_reg_in(
        ID_pipeline_reg_out), .pipeline_reg_out(EX_pipeline_reg_out) );
  MEM_stage MEM_stage_inst ( .clk(clk), .rst(n4), .pipeline_reg_in(
        EX_pipeline_reg_out), .pipeline_reg_out(MEM_pipeline_reg_out) );
  WB_stage WB_stage_inst ( .clk(clk), .rst(n4), .pipeline_reg_in(
        MEM_pipeline_reg_out), .reg_write_en(reg_write_en), .reg_write_dest(
        reg_write_dest), .reg_write_data(reg_write_data), 
        .instruction_fetch_en(instruction_fetch_en) );
  register_file register_file_inst ( .clk(clk), .rst(n4), .reg_write_en(
        reg_write_en), .reg_write_dest(reg_write_dest), .reg_write_data(
        reg_write_data), .reg_read_addr_1({n1, reg_read_addr_1[1:0]}), 
        .reg_read_data_1(reg_read_data_1), .reg_read_addr_2(reg_read_addr_2), 
        .reg_read_data_2(reg_read_data_2) );
  BUFX2 U1 ( .A(reg_read_addr_1[2]), .Y(n1) );
  INVX2 U2 ( .A(n3), .Y(n4) );
  INVX2 U3 ( .A(rst), .Y(n3) );
endmodule

